-- cineraria_core.vhd

-- Generated using ACDS version 13.0sp1 232 at 2013.10.15.04:24:49

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cineraria_core is
	port (
		clk_100mhz_clk    : in    std_logic                     := '0';             -- clk_100mhz.clk
		sys_reset_reset_n : in    std_logic                     := '0';             --  sys_reset.reset_n
		clk_40mhz_clk     : in    std_logic                     := '0';             --  clk_40mhz.clk
		sysuart_rxd       : in    std_logic                     := '0';             --    sysuart.rxd
		sysuart_txd       : out   std_logic;                                        --           .txd
		sysuart_cts_n     : in    std_logic                     := '0';             --           .cts_n
		sysuart_rts_n     : out   std_logic;                                        --           .rts_n
		sdr_addr          : out   std_logic_vector(11 downto 0);                    --        sdr.addr
		sdr_ba            : out   std_logic_vector(1 downto 0);                     --           .ba
		sdr_cas_n         : out   std_logic;                                        --           .cas_n
		sdr_cke           : out   std_logic;                                        --           .cke
		sdr_cs_n          : out   std_logic;                                        --           .cs_n
		sdr_dq            : inout std_logic_vector(15 downto 0) := (others => '0'); --           .dq
		sdr_dqm           : out   std_logic_vector(1 downto 0);                     --           .dqm
		sdr_ras_n         : out   std_logic;                                        --           .ras_n
		sdr_we_n          : out   std_logic;                                        --           .we_n
		led_export        : out   std_logic_vector(9 downto 0);                     --        led.export
		led_7seg_export   : out   std_logic_vector(31 downto 0);                    --   led_7seg.export
		psw_export        : in    std_logic_vector(2 downto 0)  := (others => '0'); --        psw.export
		dipsw_export      : in    std_logic_vector(9 downto 0)  := (others => '0'); --      dipsw.export
		spu_clk_128fs     : in    std_logic                     := '0';             --        spu.clk_128fs
		spu_DAC_BCLK      : out   std_logic;                                        --           .DAC_BCLK
		spu_DAC_LRCK      : out   std_logic;                                        --           .DAC_LRCK
		spu_DAC_DATA      : out   std_logic;                                        --           .DAC_DATA
		spu_AUD_L         : out   std_logic;                                        --           .AUD_L
		spu_AUD_R         : out   std_logic;                                        --           .AUD_R
		spu_SPDIF         : out   std_logic;                                        --           .SPDIF
		mmc_nCS           : out   std_logic;                                        --        mmc.nCS
		mmc_SCK           : out   std_logic;                                        --           .SCK
		mmc_SDO           : out   std_logic;                                        --           .SDO
		mmc_SDI           : in    std_logic                     := '0';             --           .SDI
		mmc_CD            : in    std_logic                     := '0';             --           .CD
		mmc_WP            : in    std_logic                     := '0';             --           .WP
		ps2kb_CLK         : inout std_logic                     := '0';             --      ps2kb.CLK
		ps2kb_DAT         : inout std_logic                     := '0';             --           .DAT
		gpio1_export      : inout std_logic_vector(31 downto 0) := (others => '0'); --      gpio1.export
		vga_clk           : in    std_logic                     := '0';             --        vga.clk
		vga_rout          : out   std_logic_vector(4 downto 0);                     --           .rout
		vga_gout          : out   std_logic_vector(4 downto 0);                     --           .gout
		vga_bout          : out   std_logic_vector(4 downto 0);                     --           .bout
		vga_hsync_n       : out   std_logic;                                        --           .hsync_n
		vga_vsync_n       : out   std_logic;                                        --           .vsync_n
		vga_enable        : out   std_logic;                                        --           .enable
		blcon_on          : out   std_logic;                                        --      blcon.on
		blcon_pwm         : out   std_logic                                         --           .pwm
	);
end entity cineraria_core;

architecture rtl of cineraria_core is
	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			ADDRESS_WIDTH       : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(13 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component cineraria_core_nios2_fast is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			A_ci_multi_done                       : in  std_logic                     := 'X';             -- done
			A_ci_multi_result                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_result
			A_ci_multi_a                          : out std_logic_vector(4 downto 0);                     -- multi_a
			A_ci_multi_b                          : out std_logic_vector(4 downto 0);                     -- multi_b
			A_ci_multi_c                          : out std_logic_vector(4 downto 0);                     -- multi_c
			A_ci_multi_clk_en                     : out std_logic;                                        -- clk_en
			A_ci_multi_clock                      : out std_logic;                                        -- clk
			A_ci_multi_reset                      : out std_logic;                                        -- reset
			A_ci_multi_dataa                      : out std_logic_vector(31 downto 0);                    -- multi_dataa
			A_ci_multi_datab                      : out std_logic_vector(31 downto 0);                    -- multi_datab
			A_ci_multi_n                          : out std_logic_vector(7 downto 0);                     -- multi_n
			A_ci_multi_readra                     : out std_logic;                                        -- multi_readra
			A_ci_multi_readrb                     : out std_logic;                                        -- multi_readrb
			A_ci_multi_start                      : out std_logic;                                        -- start
			A_ci_multi_writerc                    : out std_logic                                         -- multi_writerc
		);
	end component cineraria_core_nios2_fast;

	component fpoint_wrapper is
		generic (
			useDivider : integer := 0
		);
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			clk_en : in  std_logic                     := 'X';             -- clk_en
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			n      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- n
			reset  : in  std_logic                     := 'X';             -- reset
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component fpoint_wrapper;

	component cineraria_core_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component cineraria_core_jtag_uart;

	component cineraria_core_sysuart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			cts_n         : in  std_logic                     := 'X';             -- export
			rts_n         : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component cineraria_core_sysuart;

	component cineraria_core_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component cineraria_core_sdram;

	component cineraria_core_ipl_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component cineraria_core_ipl_memory;

	component cineraria_core_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component cineraria_core_sysid;

	component cineraria_core_systimer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component cineraria_core_systimer;

	component cineraria_core_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component cineraria_core_led;

	component cineraria_core_led_7seg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component cineraria_core_led_7seg;

	component cineraria_core_psw is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component cineraria_core_psw;

	component cineraria_core_dipsw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component cineraria_core_dipsw;

	component pixelsimd is
		port (
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			result : out std_logic_vector(31 downto 0);                    -- result
			clk    : in  std_logic                     := 'X';             -- clk
			clk_en : in  std_logic                     := 'X';             -- clk_en
			reset  : in  std_logic                     := 'X';             -- reset
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			n      : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- n
		);
	end component pixelsimd;

	component avalonif_spu is
		port (
			csi_global_clock     : in  std_logic                     := 'X';             -- clk
			csi_global_reset     : in  std_logic                     := 'X';             -- reset
			csi_m1_clock         : in  std_logic                     := 'X';             -- clk
			avm_m1_address       : out std_logic_vector(24 downto 0);                    -- address
			avm_m1_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			avm_m1_read          : out std_logic;                                        -- read
			avm_m1_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avm_m1_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avm_m1_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avs_s1_address       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			avs_s1_chipselect    : in  std_logic                     := 'X';             -- chipselect
			avs_s1_read          : in  std_logic                     := 'X';             -- read
			avs_s1_write         : in  std_logic                     := 'X';             -- write
			avs_s1_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s1_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s1_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s1_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s1_irq           : out std_logic;                                        -- irq
			clk_128fs            : in  std_logic                     := 'X';             -- export
			DAC_BCLK             : out std_logic;                                        -- export
			DAC_LRCK             : out std_logic;                                        -- export
			DAC_DATA             : out std_logic;                                        -- export
			AUD_L                : out std_logic;                                        -- export
			AUD_R                : out std_logic;                                        -- export
			SPDIF                : out std_logic                                         -- export
		);
	end component avalonif_spu;

	component avalonif_mmcdma is
		generic (
			SYSTEMCLOCKINFO : integer := 0
		);
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			chipselect : in  std_logic                     := 'X';             -- chipselect
			address    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			read       : in  std_logic                     := 'X';             -- read
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			MMC_nCS    : out std_logic;                                        -- export
			MMC_SCK    : out std_logic;                                        -- export
			MMC_SDO    : out std_logic;                                        -- export
			MMC_SDI    : in  std_logic                     := 'X';             -- export
			MMC_CD     : in  std_logic                     := 'X';             -- export
			MMC_WP     : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component avalonif_mmcdma;

	component ps2_component is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X';             -- export
			irq         : out   std_logic                                         -- irq
		);
	end component ps2_component;

	component cineraria_core_gpio1 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component cineraria_core_gpio1;

	component vga_component is
		generic (
			LINEOFFSETBYTES : integer := 2048;
			H_TOTAL         : integer := 800;
			H_SYNC          : integer := 96;
			H_BACKP         : integer := 48;
			H_ACTIVE        : integer := 640;
			V_TOTAL         : integer := 525;
			V_SYNC          : integer := 2;
			V_BACKP         : integer := 33;
			V_ACTIVE        : integer := 480
		);
		port (
			video_clk            : in  std_logic                     := 'X';             -- export
			video_rout           : out std_logic_vector(4 downto 0);                     -- export
			video_gout           : out std_logic_vector(4 downto 0);                     -- export
			video_bout           : out std_logic_vector(4 downto 0);                     -- export
			video_hsync_n        : out std_logic;                                        -- export
			video_vsync_n        : out std_logic;                                        -- export
			video_enable         : out std_logic;                                        -- export
			avm_m1_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_m1_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_m1_burstcount    : out std_logic_vector(9 downto 0);                     -- burstcount
			avm_m1_read          : out std_logic;                                        -- read
			avm_m1_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_m1_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avs_s1_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_s1_read          : in  std_logic                     := 'X';             -- read
			avs_s1_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s1_write         : in  std_logic                     := 'X';             -- write
			avs_s1_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq_s1               : out std_logic;                                        -- irq
			s1_clk               : in  std_logic                     := 'X';             -- clk
			m1_clk               : in  std_logic                     := 'X';             -- clk
			g_reset              : in  std_logic                     := 'X'              -- reset
		);
	end component vga_component;

	component backlight_control is
		port (
			reset         : in  std_logic                     := 'X';             -- reset
			clk           : in  std_logic                     := 'X';             -- clk
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			backlight_on  : out std_logic;                                        -- export
			backlight_pwm : out std_logic                                         -- export
		);
	end component backlight_control;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_result         : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_multi_clk      : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset    : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken    : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_start    : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done     : out std_logic;                                        -- done
			ci_slave_multi_dataa    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result   : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra   : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb   : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc  : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_c
			comb_ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_clk     : out std_logic;                                        -- clk
			multi_ci_master_reset   : out std_logic;                                        -- reset
			multi_ci_master_clken   : out std_logic;                                        -- clk_en
			multi_ci_master_start   : out std_logic;                                        -- start
			multi_ci_master_done    : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa   : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab   : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n       : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra  : out std_logic;                                        -- readra
			multi_ci_master_readrb  : out std_logic;                                        -- readrb
			multi_ci_master_writerc : out std_logic;                                        -- writerc
			multi_ci_master_a       : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b       : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c       : out std_logic_vector(4 downto 0);                     -- c
			ci_slave_dataa          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_n              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra         : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb         : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc        : in  std_logic                     := 'X';             -- writerc
			ci_slave_a              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus        : in  std_logic                     := 'X';             -- estatus
			comb_ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab    : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_n        : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra   : out std_logic;                                        -- readra
			comb_ci_master_readrb   : out std_logic;                                        -- readrb
			comb_ci_master_writerc  : out std_logic;                                        -- writerc
			comb_ci_master_a        : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b        : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c        : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus  : out std_logic                                         -- estatus
		);
	end component altera_customins_master_translator;

	component cineraria_core_nios2_fast_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic;                                        -- done
			ci_master0_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra   : out std_logic;                                        -- readra
			ci_master0_readrb   : out std_logic;                                        -- readrb
			ci_master0_writerc  : out std_logic;                                        -- writerc
			ci_master0_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus  : out std_logic;                                        -- estatus
			ci_master0_clk      : out std_logic;                                        -- clk
			ci_master0_reset    : out std_logic;                                        -- reset
			ci_master0_clken    : out std_logic;                                        -- clk_en
			ci_master0_start    : out std_logic;                                        -- start
			ci_master0_done     : in  std_logic                     := 'X';             -- done
			ci_master1_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master1_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master1_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master1_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master1_readra   : out std_logic;                                        -- readra
			ci_master1_readrb   : out std_logic;                                        -- readrb
			ci_master1_writerc  : out std_logic;                                        -- writerc
			ci_master1_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master1_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master1_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master1_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master1_estatus  : out std_logic;                                        -- estatus
			ci_master1_clk      : out std_logic;                                        -- clk
			ci_master1_reset    : out std_logic;                                        -- reset
			ci_master1_clken    : out std_logic;                                        -- clk_en
			ci_master1_start    : out std_logic;                                        -- start
			ci_master1_done     : in  std_logic                     := 'X'              -- done
		);
	end component cineraria_core_nios2_fast_custom_instruction_master_multi_xconnect;

	component cineraria_core_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(114 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_addr_router;

	component cineraria_core_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(114 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_addr_router_001;

	component cineraria_core_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(96 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_addr_router_002;

	component cineraria_core_addr_router_003 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(114 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_addr_router_003;

	component cineraria_core_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(114 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_id_router;

	component cineraria_core_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(96 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_id_router_002;

	component cineraria_core_id_router_003 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(114 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_id_router_003;

	component cineraria_core_addr_router_004 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(86 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_addr_router_004;

	component cineraria_core_id_router_004 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(86 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_id_router_004;

	component cineraria_core_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(114 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(114 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(114 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_cmd_xbar_demux;

	component cineraria_core_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(114 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(114 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(114 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(114 downto 0);                    -- data
			src3_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_cmd_xbar_demux_001;

	component cineraria_core_cmd_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(96 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_cmd_xbar_demux_002;

	component cineraria_core_cmd_xbar_demux_003 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(114 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_cmd_xbar_demux_003;

	component cineraria_core_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(114 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component cineraria_core_cmd_xbar_mux;

	component cineraria_core_cmd_xbar_mux_002 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(96 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component cineraria_core_cmd_xbar_mux_002;

	component cineraria_core_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(114 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(114 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component cineraria_core_rsp_xbar_demux;

	component cineraria_core_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(96 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(96 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(96 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(96 downto 0);                    -- data
			src3_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_rsp_xbar_demux_002;

	component cineraria_core_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(114 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component cineraria_core_rsp_xbar_mux;

	component cineraria_core_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(114 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component cineraria_core_rsp_xbar_mux_001;

	component cineraria_core_cmd_xbar_demux_004 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(13 downto 0) := (others => 'X'); -- data
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(86 downto 0);                    -- data
			src0_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(86 downto 0);                    -- data
			src1_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(86 downto 0);                    -- data
			src2_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(86 downto 0);                    -- data
			src3_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(86 downto 0);                    -- data
			src4_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(86 downto 0);                    -- data
			src5_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(86 downto 0);                    -- data
			src6_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(86 downto 0);                    -- data
			src7_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(86 downto 0);                    -- data
			src8_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(86 downto 0);                    -- data
			src9_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(86 downto 0);                    -- data
			src10_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(86 downto 0);                    -- data
			src11_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(86 downto 0);                    -- data
			src12_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(86 downto 0);                    -- data
			src13_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_cmd_xbar_demux_004;

	component cineraria_core_rsp_xbar_demux_004 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(86 downto 0);                    -- data
			src0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cineraria_core_rsp_xbar_demux_004;

	component cineraria_core_rsp_xbar_mux_004 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(86 downto 0);                    -- data
			src_channel          : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component cineraria_core_rsp_xbar_mux_004;

	component cineraria_core_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component cineraria_core_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component cineraria_core_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(114 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(114 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(3 downto 0)                       -- data
		);
	end component cineraria_core_limiter;

	component cineraria_core_limiter_002 is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(86 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(86 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(13 downto 0)                     -- data
		);
	end component cineraria_core_limiter_002;

	component cineraria_core_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(96 downto 0);                     -- data
			out_channel          : out std_logic_vector(3 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component cineraria_core_width_adapter;

	component cineraria_core_width_adapter_003 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(96 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(114 downto 0);                    -- data
			out_channel          : out std_logic_vector(3 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component cineraria_core_width_adapter_003;

	component cineraria_core_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                      := 'X';             -- clk
			reset                 : in  std_logic                      := 'X';             -- reset
			sink0_valid           : in  std_logic                      := 'X';             -- valid
			sink0_data            : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                         -- ready
			source0_valid         : out std_logic;                                         -- valid
			source0_data          : out std_logic_vector(114 downto 0);                    -- data
			source0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			source0_startofpacket : out std_logic;                                         -- startofpacket
			source0_endofpacket   : out std_logic;                                         -- endofpacket
			source0_ready         : in  std_logic                      := 'X'              -- ready
		);
	end component cineraria_core_burst_adapter;

	component cineraria_core_burst_adapter_002 is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(96 downto 0);                    -- data
			source0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component cineraria_core_burst_adapter_002;

	component cineraria_core_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component cineraria_core_rst_controller;

	component cineraria_core_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component cineraria_core_rst_controller_001;

	component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(115 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(115 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(33 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(97 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(87 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(87 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(114 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(115 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(115 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(96 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(97 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent;

	component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(13 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(86 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(87 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(87 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent;

	component cineraria_core_nios2_fast_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(5 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_nios2_fast_instruction_master_translator;

	component cineraria_core_nios2_fast_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(5 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_nios2_fast_data_master_translator;

	component cineraria_core_spu_m1_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(3 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(15 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_byteenable            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_spu_m1_translator;

	component cineraria_core_vga_m1_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(11 downto 0);                    -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- burstcount
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_vga_m1_translator;

	component cineraria_core_peripherals_bridge_m0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(13 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_peripherals_bridge_m0_translator;

	component cineraria_core_nios2_fast_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_nios2_fast_jtag_debug_module_translator;

	component cineraria_core_ipl_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(10 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_ipl_memory_s1_translator;

	component cineraria_core_sdram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_sdram_s1_translator;

	component cineraria_core_peripherals_bridge_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(13 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_peripherals_bridge_s0_translator;

	component cineraria_core_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_jtag_uart_avalon_jtag_slave_translator;

	component cineraria_core_sysuart_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_chipselect            : out std_logic;                                        -- chipselect
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_sysuart_s1_translator;

	component cineraria_core_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_sysid_control_slave_translator;

	component cineraria_core_systimer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_systimer_s1_translator;

	component cineraria_core_led_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_led_s1_translator;

	component cineraria_core_dipsw_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_dipsw_s1_translator;

	component cineraria_core_spu_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_spu_s1_translator;

	component cineraria_core_mmcdma_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_mmcdma_s1_translator;

	component cineraria_core_ps2_keyboard_avalon_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_ps2_keyboard_avalon_slave_translator;

	component cineraria_core_vga_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_vga_s1_translator;

	component cineraria_core_blcon_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cineraria_core_blcon_s1_translator;

	component cineraria_core_nios2_fast_instruction_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(114 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component cineraria_core_nios2_fast_instruction_master_translator_avalon_universal_master_0_agent;

	component cineraria_core_spu_m1_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(96 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_spu_m1_translator_avalon_universal_master_0_agent;

	component cineraria_core_vga_m1_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(114 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(114 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component cineraria_core_vga_m1_translator_avalon_universal_master_0_agent;

	component cineraria_core_peripherals_bridge_m0_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(86 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component cineraria_core_peripherals_bridge_m0_translator_avalon_universal_master_0_agent;

	component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator0 is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result    : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra    : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb    : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc   : in  std_logic                     := 'X';             -- writerc
			ci_slave_a         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus   : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk       : in  std_logic                     := 'X';             -- clk
			ci_slave_clken     : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset     : in  std_logic                     := 'X';             -- reset
			ci_slave_start     : in  std_logic                     := 'X';             -- start
			ci_slave_done      : out std_logic;                                        -- done
			ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n        : out std_logic_vector(1 downto 0);                     -- n
			ci_master_clk      : out std_logic;                                        -- clk
			ci_master_clken    : out std_logic;                                        -- clk_en
			ci_master_reset    : out std_logic;                                        -- reset
			ci_master_start    : out std_logic;                                        -- start
			ci_master_done     : in  std_logic                     := 'X';             -- done
			ci_master_readra   : out std_logic;                                        -- readra
			ci_master_readrb   : out std_logic;                                        -- readrb
			ci_master_writerc  : out std_logic;                                        -- writerc
			ci_master_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus  : out std_logic                                         -- estatus
		);
	end component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator0;

	component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator1 is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result    : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra    : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb    : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc   : in  std_logic                     := 'X';             -- writerc
			ci_slave_a         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus   : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk       : in  std_logic                     := 'X';             -- clk
			ci_slave_clken     : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset     : in  std_logic                     := 'X';             -- reset
			ci_slave_start     : in  std_logic                     := 'X';             -- start
			ci_slave_done      : out std_logic;                                        -- done
			ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n        : out std_logic_vector(2 downto 0);                     -- n
			ci_master_clk      : out std_logic;                                        -- clk
			ci_master_clken    : out std_logic;                                        -- clk_en
			ci_master_reset    : out std_logic;                                        -- reset
			ci_master_start    : out std_logic;                                        -- start
			ci_master_done     : in  std_logic                     := 'X';             -- done
			ci_master_readra   : out std_logic;                                        -- readra
			ci_master_readrb   : out std_logic;                                        -- readrb
			ci_master_writerc  : out std_logic;                                        -- writerc
			ci_master_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus  : out std_logic                                         -- estatus
		);
	end component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator1;

	signal nios2_fast_custom_instruction_master_multi_readra                                                 : std_logic;                      -- nios2_fast:A_ci_multi_readra -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_readra
	signal nios2_fast_custom_instruction_master_multi_n                                                      : std_logic_vector(7 downto 0);   -- nios2_fast:A_ci_multi_n -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_n
	signal nios2_fast_custom_instruction_master_multi_readrb                                                 : std_logic;                      -- nios2_fast:A_ci_multi_readrb -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_readrb
	signal nios2_fast_custom_instruction_master_done                                                         : std_logic;                      -- nios2_fast_custom_instruction_master_translator:ci_slave_multi_done -> nios2_fast:A_ci_multi_done
	signal nios2_fast_custom_instruction_master_clk_en                                                       : std_logic;                      -- nios2_fast:A_ci_multi_clk_en -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_clken
	signal nios2_fast_custom_instruction_master_multi_writerc                                                : std_logic;                      -- nios2_fast:A_ci_multi_writerc -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_writerc
	signal nios2_fast_custom_instruction_master_multi_result                                                 : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_translator:ci_slave_multi_result -> nios2_fast:A_ci_multi_result
	signal nios2_fast_custom_instruction_master_clk                                                          : std_logic;                      -- nios2_fast:A_ci_multi_clock -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_clk
	signal nios2_fast_custom_instruction_master_multi_c                                                      : std_logic_vector(4 downto 0);   -- nios2_fast:A_ci_multi_c -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_c
	signal nios2_fast_custom_instruction_master_multi_b                                                      : std_logic_vector(4 downto 0);   -- nios2_fast:A_ci_multi_b -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_b
	signal nios2_fast_custom_instruction_master_multi_a                                                      : std_logic_vector(4 downto 0);   -- nios2_fast:A_ci_multi_a -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_a
	signal nios2_fast_custom_instruction_master_multi_dataa                                                  : std_logic_vector(31 downto 0);  -- nios2_fast:A_ci_multi_dataa -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_dataa
	signal nios2_fast_custom_instruction_master_start                                                        : std_logic;                      -- nios2_fast:A_ci_multi_start -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_start
	signal nios2_fast_custom_instruction_master_multi_datab                                                  : std_logic_vector(31 downto 0);  -- nios2_fast:A_ci_multi_datab -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_datab
	signal nios2_fast_custom_instruction_master_reset                                                        : std_logic;                      -- nios2_fast:A_ci_multi_reset -> nios2_fast_custom_instruction_master_translator:ci_slave_multi_reset
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_result                            : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_fast_custom_instruction_master_translator:multi_ci_master_result
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_b                                 : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_translator:multi_ci_master_b -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_b
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_c                                 : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_translator:multi_ci_master_c -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_c
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en                            : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_clken -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_done                              : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_fast_custom_instruction_master_translator:multi_ci_master_done
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_a                                 : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_translator:multi_ci_master_a -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_a
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_n                                 : std_logic_vector(7 downto 0);   -- nios2_fast_custom_instruction_master_translator:multi_ci_master_n -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_n
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc                           : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_clk                               : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_clk -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_start                             : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_start -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_start
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa                             : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_readra                            : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_readra -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_reset                             : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_reset -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_datab                             : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_translator:multi_ci_master_datab -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb                            : std_logic;                      -- nios2_fast_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_fast_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result                             : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_result
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done                               : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_done
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n                                  : std_logic_vector(7 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc                            : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending                           : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk                                : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start                              : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa                              : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset                              : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab                              : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus                            : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result                     : std_logic_vector(31 downto 0);  -- nios_custom_instr_fpoint:result -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start                      : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_fpoint:start
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa                      : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_fpoint:dataa
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done                       : std_logic;                      -- nios_custom_instr_fpoint:done -> nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en                     : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_fpoint:clk_en
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n                          : std_logic_vector(1 downto 0);   -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_fpoint:n
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset                      : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_fpoint:reset
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab                      : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_fpoint:datab
	signal nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk                        : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_fpoint:clk
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result                             : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_result
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_b
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_c
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done                               : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_done
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a                                  : std_logic_vector(4 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_a
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n                                  : std_logic_vector(7 downto 0);   -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_n
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc                            : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending                           : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk                                : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start                              : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_start
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa                              : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset                              : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab                              : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb                             : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	signal nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus                            : std_logic;                      -- nios2_fast_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result                     : std_logic_vector(31 downto 0);  -- nios_custom_instr_pixelsimd:result -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_result
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start                      : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_start -> nios_custom_instr_pixelsimd:start
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa                      : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> nios_custom_instr_pixelsimd:dataa
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done                       : std_logic;                      -- nios_custom_instr_pixelsimd:done -> nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_done
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en                     : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_clken -> nios_custom_instr_pixelsimd:clk_en
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n                          : std_logic_vector(2 downto 0);   -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_n -> nios_custom_instr_pixelsimd:n
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset                      : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_reset -> nios_custom_instr_pixelsimd:reset
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab                      : std_logic_vector(31 downto 0);  -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_datab -> nios_custom_instr_pixelsimd:datab
	signal nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk                        : std_logic;                      -- nios2_fast_custom_instruction_master_multi_slave_translator1:ci_master_clk -> nios_custom_instr_pixelsimd:clk
	signal nios2_fast_instruction_master_burstcount                                                          : std_logic_vector(3 downto 0);   -- nios2_fast:i_burstcount -> nios2_fast_instruction_master_translator:av_burstcount
	signal nios2_fast_instruction_master_waitrequest                                                         : std_logic;                      -- nios2_fast_instruction_master_translator:av_waitrequest -> nios2_fast:i_waitrequest
	signal nios2_fast_instruction_master_address                                                             : std_logic_vector(27 downto 0);  -- nios2_fast:i_address -> nios2_fast_instruction_master_translator:av_address
	signal nios2_fast_instruction_master_read                                                                : std_logic;                      -- nios2_fast:i_read -> nios2_fast_instruction_master_translator:av_read
	signal nios2_fast_instruction_master_readdata                                                            : std_logic_vector(31 downto 0);  -- nios2_fast_instruction_master_translator:av_readdata -> nios2_fast:i_readdata
	signal nios2_fast_instruction_master_readdatavalid                                                       : std_logic;                      -- nios2_fast_instruction_master_translator:av_readdatavalid -> nios2_fast:i_readdatavalid
	signal nios2_fast_data_master_burstcount                                                                 : std_logic_vector(3 downto 0);   -- nios2_fast:d_burstcount -> nios2_fast_data_master_translator:av_burstcount
	signal nios2_fast_data_master_waitrequest                                                                : std_logic;                      -- nios2_fast_data_master_translator:av_waitrequest -> nios2_fast:d_waitrequest
	signal nios2_fast_data_master_writedata                                                                  : std_logic_vector(31 downto 0);  -- nios2_fast:d_writedata -> nios2_fast_data_master_translator:av_writedata
	signal nios2_fast_data_master_address                                                                    : std_logic_vector(28 downto 0);  -- nios2_fast:d_address -> nios2_fast_data_master_translator:av_address
	signal nios2_fast_data_master_write                                                                      : std_logic;                      -- nios2_fast:d_write -> nios2_fast_data_master_translator:av_write
	signal nios2_fast_data_master_read                                                                       : std_logic;                      -- nios2_fast:d_read -> nios2_fast_data_master_translator:av_read
	signal nios2_fast_data_master_readdata                                                                   : std_logic_vector(31 downto 0);  -- nios2_fast_data_master_translator:av_readdata -> nios2_fast:d_readdata
	signal nios2_fast_data_master_debugaccess                                                                : std_logic;                      -- nios2_fast:jtag_debug_module_debugaccess_to_roms -> nios2_fast_data_master_translator:av_debugaccess
	signal nios2_fast_data_master_readdatavalid                                                              : std_logic;                      -- nios2_fast_data_master_translator:av_readdatavalid -> nios2_fast:d_readdatavalid
	signal nios2_fast_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);   -- nios2_fast:d_byteenable -> nios2_fast_data_master_translator:av_byteenable
	signal spu_m1_waitrequest                                                                                : std_logic;                      -- spu_m1_translator:av_waitrequest -> spu:avm_m1_waitrequest
	signal spu_m1_burstcount                                                                                 : std_logic_vector(2 downto 0);   -- spu:avm_m1_burstcount -> spu_m1_translator:av_burstcount
	signal spu_m1_address                                                                                    : std_logic_vector(24 downto 0);  -- spu:avm_m1_address -> spu_m1_translator:av_address
	signal spu_m1_read                                                                                       : std_logic;                      -- spu:avm_m1_read -> spu_m1_translator:av_read
	signal spu_m1_readdata                                                                                   : std_logic_vector(15 downto 0);  -- spu_m1_translator:av_readdata -> spu:avm_m1_readdata
	signal spu_m1_readdatavalid                                                                              : std_logic;                      -- spu_m1_translator:av_readdatavalid -> spu:avm_m1_readdatavalid
	signal vga_m1_burstcount                                                                                 : std_logic_vector(9 downto 0);   -- vga:avm_m1_burstcount -> vga_m1_translator:av_burstcount
	signal vga_m1_waitrequest                                                                                : std_logic;                      -- vga_m1_translator:av_waitrequest -> vga:avm_m1_waitrequest
	signal vga_m1_address                                                                                    : std_logic_vector(31 downto 0);  -- vga:avm_m1_address -> vga_m1_translator:av_address
	signal vga_m1_read                                                                                       : std_logic;                      -- vga:avm_m1_read -> vga_m1_translator:av_read
	signal vga_m1_readdata                                                                                   : std_logic_vector(31 downto 0);  -- vga_m1_translator:av_readdata -> vga:avm_m1_readdata
	signal vga_m1_readdatavalid                                                                              : std_logic;                      -- vga_m1_translator:av_readdatavalid -> vga:avm_m1_readdatavalid
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- nios2_fast:jtag_debug_module_waitrequest -> nios2_fast_jtag_debug_module_translator:av_waitrequest
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_fast_jtag_debug_module_translator:av_writedata -> nios2_fast:jtag_debug_module_writedata
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);   -- nios2_fast_jtag_debug_module_translator:av_address -> nios2_fast:jtag_debug_module_address
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- nios2_fast_jtag_debug_module_translator:av_write -> nios2_fast:jtag_debug_module_write
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- nios2_fast_jtag_debug_module_translator:av_read -> nios2_fast:jtag_debug_module_read
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_fast:jtag_debug_module_readdata -> nios2_fast_jtag_debug_module_translator:av_readdata
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                      -- nios2_fast_jtag_debug_module_translator:av_debugaccess -> nios2_fast:jtag_debug_module_debugaccess
	signal nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_fast_jtag_debug_module_translator:av_byteenable -> nios2_fast:jtag_debug_module_byteenable
	signal ipl_memory_s1_translator_avalon_anti_slave_0_writedata                                            : std_logic_vector(31 downto 0);  -- ipl_memory_s1_translator:av_writedata -> ipl_memory:writedata
	signal ipl_memory_s1_translator_avalon_anti_slave_0_address                                              : std_logic_vector(10 downto 0);  -- ipl_memory_s1_translator:av_address -> ipl_memory:address
	signal ipl_memory_s1_translator_avalon_anti_slave_0_chipselect                                           : std_logic;                      -- ipl_memory_s1_translator:av_chipselect -> ipl_memory:chipselect
	signal ipl_memory_s1_translator_avalon_anti_slave_0_clken                                                : std_logic;                      -- ipl_memory_s1_translator:av_clken -> ipl_memory:clken
	signal ipl_memory_s1_translator_avalon_anti_slave_0_write                                                : std_logic;                      -- ipl_memory_s1_translator:av_write -> ipl_memory:write
	signal ipl_memory_s1_translator_avalon_anti_slave_0_readdata                                             : std_logic_vector(31 downto 0);  -- ipl_memory:readdata -> ipl_memory_s1_translator:av_readdata
	signal ipl_memory_s1_translator_avalon_anti_slave_0_byteenable                                           : std_logic_vector(3 downto 0);   -- ipl_memory_s1_translator:av_byteenable -> ipl_memory:byteenable
	signal sdram_s1_translator_avalon_anti_slave_0_waitrequest                                               : std_logic;                      -- sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	signal sdram_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0);  -- sdram_s1_translator:av_writedata -> sdram:az_data
	signal sdram_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(21 downto 0);  -- sdram_s1_translator:av_address -> sdram:az_addr
	signal sdram_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- sdram_s1_translator:av_chipselect -> sdram:az_cs
	signal sdram_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- sdram_s1_translator:av_write -> sdram_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_s1_translator_avalon_anti_slave_0_read                                                      : std_logic;                      -- sdram_s1_translator:av_read -> sdram_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0);  -- sdram:za_data -> sdram_s1_translator:av_readdata
	signal sdram_s1_translator_avalon_anti_slave_0_readdatavalid                                             : std_logic;                      -- sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable                                                : std_logic_vector(1 downto 0);   -- sdram_s1_translator:av_byteenable -> sdram_s1_translator_avalon_anti_slave_0_byteenable:in
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_waitrequest                                  : std_logic;                      -- peripherals_bridge:s0_waitrequest -> peripherals_bridge_s0_translator:av_waitrequest
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_burstcount                                   : std_logic_vector(0 downto 0);   -- peripherals_bridge_s0_translator:av_burstcount -> peripherals_bridge:s0_burstcount
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- peripherals_bridge_s0_translator:av_writedata -> peripherals_bridge:s0_writedata
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_address                                      : std_logic_vector(13 downto 0);  -- peripherals_bridge_s0_translator:av_address -> peripherals_bridge:s0_address
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- peripherals_bridge_s0_translator:av_write -> peripherals_bridge:s0_write
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_read                                         : std_logic;                      -- peripherals_bridge_s0_translator:av_read -> peripherals_bridge:s0_read
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- peripherals_bridge:s0_readdata -> peripherals_bridge_s0_translator:av_readdata
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_debugaccess                                  : std_logic;                      -- peripherals_bridge_s0_translator:av_debugaccess -> peripherals_bridge:s0_debugaccess
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_readdatavalid                                : std_logic;                      -- peripherals_bridge:s0_readdatavalid -> peripherals_bridge_s0_translator:av_readdatavalid
	signal peripherals_bridge_s0_translator_avalon_anti_slave_0_byteenable                                   : std_logic_vector(3 downto 0);   -- peripherals_bridge_s0_translator:av_byteenable -> peripherals_bridge:s0_byteenable
	signal peripherals_bridge_m0_burstcount                                                                  : std_logic_vector(0 downto 0);   -- peripherals_bridge:m0_burstcount -> peripherals_bridge_m0_translator:av_burstcount
	signal peripherals_bridge_m0_waitrequest                                                                 : std_logic;                      -- peripherals_bridge_m0_translator:av_waitrequest -> peripherals_bridge:m0_waitrequest
	signal peripherals_bridge_m0_address                                                                     : std_logic_vector(13 downto 0);  -- peripherals_bridge:m0_address -> peripherals_bridge_m0_translator:av_address
	signal peripherals_bridge_m0_writedata                                                                   : std_logic_vector(31 downto 0);  -- peripherals_bridge:m0_writedata -> peripherals_bridge_m0_translator:av_writedata
	signal peripherals_bridge_m0_write                                                                       : std_logic;                      -- peripherals_bridge:m0_write -> peripherals_bridge_m0_translator:av_write
	signal peripherals_bridge_m0_read                                                                        : std_logic;                      -- peripherals_bridge:m0_read -> peripherals_bridge_m0_translator:av_read
	signal peripherals_bridge_m0_readdata                                                                    : std_logic_vector(31 downto 0);  -- peripherals_bridge_m0_translator:av_readdata -> peripherals_bridge:m0_readdata
	signal peripherals_bridge_m0_debugaccess                                                                 : std_logic;                      -- peripherals_bridge:m0_debugaccess -> peripherals_bridge_m0_translator:av_debugaccess
	signal peripherals_bridge_m0_byteenable                                                                  : std_logic_vector(3 downto 0);   -- peripherals_bridge:m0_byteenable -> peripherals_bridge_m0_translator:av_byteenable
	signal peripherals_bridge_m0_readdatavalid                                                               : std_logic;                      -- peripherals_bridge_m0_translator:av_readdatavalid -> peripherals_bridge:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                      -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);   -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal sysuart_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(15 downto 0);  -- sysuart_s1_translator:av_writedata -> sysuart:writedata
	signal sysuart_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(2 downto 0);   -- sysuart_s1_translator:av_address -> sysuart:address
	signal sysuart_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                      -- sysuart_s1_translator:av_chipselect -> sysuart:chipselect
	signal sysuart_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                      -- sysuart_s1_translator:av_write -> sysuart_s1_translator_avalon_anti_slave_0_write:in
	signal sysuart_s1_translator_avalon_anti_slave_0_read                                                    : std_logic;                      -- sysuart_s1_translator:av_read -> sysuart_s1_translator_avalon_anti_slave_0_read:in
	signal sysuart_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(15 downto 0);  -- sysuart:readdata -> sysuart_s1_translator:av_readdata
	signal sysuart_s1_translator_avalon_anti_slave_0_begintransfer                                           : std_logic;                      -- sysuart_s1_translator:av_begintransfer -> sysuart:begintransfer
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                        : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal systimer_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(15 downto 0);  -- systimer_s1_translator:av_writedata -> systimer:writedata
	signal systimer_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(2 downto 0);   -- systimer_s1_translator:av_address -> systimer:address
	signal systimer_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                      -- systimer_s1_translator:av_chipselect -> systimer:chipselect
	signal systimer_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                      -- systimer_s1_translator:av_write -> systimer_s1_translator_avalon_anti_slave_0_write:in
	signal systimer_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(15 downto 0);  -- systimer:readdata -> systimer_s1_translator:av_readdata
	signal led_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- led_s1_translator:av_writedata -> led:writedata
	signal led_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- led_s1_translator:av_address -> led:address
	signal led_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- led_s1_translator:av_chipselect -> led:chipselect
	signal led_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- led_s1_translator:av_write -> led_s1_translator_avalon_anti_slave_0_write:in
	signal led_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- led:readdata -> led_s1_translator:av_readdata
	signal led_7seg_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0);  -- led_7seg_s1_translator:av_writedata -> led_7seg:writedata
	signal led_7seg_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(1 downto 0);   -- led_7seg_s1_translator:av_address -> led_7seg:address
	signal led_7seg_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                      -- led_7seg_s1_translator:av_chipselect -> led_7seg:chipselect
	signal led_7seg_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                      -- led_7seg_s1_translator:av_write -> led_7seg_s1_translator_avalon_anti_slave_0_write:in
	signal led_7seg_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0);  -- led_7seg:readdata -> led_7seg_s1_translator:av_readdata
	signal psw_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- psw_s1_translator:av_writedata -> psw:writedata
	signal psw_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- psw_s1_translator:av_address -> psw:address
	signal psw_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- psw_s1_translator:av_chipselect -> psw:chipselect
	signal psw_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- psw_s1_translator:av_write -> psw_s1_translator_avalon_anti_slave_0_write:in
	signal psw_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- psw:readdata -> psw_s1_translator:av_readdata
	signal dipsw_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);   -- dipsw_s1_translator:av_address -> dipsw:address
	signal dipsw_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- dipsw:readdata -> dipsw_s1_translator:av_readdata
	signal spu_s1_translator_avalon_anti_slave_0_waitrequest                                                 : std_logic;                      -- spu:avs_s1_waitrequest -> spu_s1_translator:av_waitrequest
	signal spu_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- spu_s1_translator:av_writedata -> spu:avs_s1_writedata
	signal spu_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(8 downto 0);   -- spu_s1_translator:av_address -> spu:avs_s1_address
	signal spu_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- spu_s1_translator:av_chipselect -> spu:avs_s1_chipselect
	signal spu_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- spu_s1_translator:av_write -> spu:avs_s1_write
	signal spu_s1_translator_avalon_anti_slave_0_read                                                        : std_logic;                      -- spu_s1_translator:av_read -> spu:avs_s1_read
	signal spu_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- spu:avs_s1_readdata -> spu_s1_translator:av_readdata
	signal spu_s1_translator_avalon_anti_slave_0_byteenable                                                  : std_logic_vector(3 downto 0);   -- spu_s1_translator:av_byteenable -> spu:avs_s1_byteenable
	signal mmcdma_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0);  -- mmcdma_s1_translator:av_writedata -> mmcdma:writedata
	signal mmcdma_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(7 downto 0);   -- mmcdma_s1_translator:av_address -> mmcdma:address
	signal mmcdma_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                      -- mmcdma_s1_translator:av_chipselect -> mmcdma:chipselect
	signal mmcdma_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                      -- mmcdma_s1_translator:av_write -> mmcdma:write
	signal mmcdma_s1_translator_avalon_anti_slave_0_read                                                     : std_logic;                      -- mmcdma_s1_translator:av_read -> mmcdma:read
	signal mmcdma_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0);  -- mmcdma:readdata -> mmcdma_s1_translator:av_readdata
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_waitrequest                              : std_logic;                      -- ps2_keyboard:waitrequest -> ps2_keyboard_avalon_slave_translator:av_waitrequest
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- ps2_keyboard_avalon_slave_translator:av_writedata -> ps2_keyboard:writedata
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_address                                  : std_logic_vector(0 downto 0);   -- ps2_keyboard_avalon_slave_translator:av_address -> ps2_keyboard:address
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- ps2_keyboard_avalon_slave_translator:av_chipselect -> ps2_keyboard:chipselect
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- ps2_keyboard_avalon_slave_translator:av_write -> ps2_keyboard:write
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_read                                     : std_logic;                      -- ps2_keyboard_avalon_slave_translator:av_read -> ps2_keyboard:read
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- ps2_keyboard:readdata -> ps2_keyboard_avalon_slave_translator:av_readdata
	signal ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);   -- ps2_keyboard_avalon_slave_translator:av_byteenable -> ps2_keyboard:byteenable
	signal gpio1_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- gpio1_s1_translator:av_writedata -> gpio1:writedata
	signal gpio1_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);   -- gpio1_s1_translator:av_address -> gpio1:address
	signal gpio1_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- gpio1_s1_translator:av_chipselect -> gpio1:chipselect
	signal gpio1_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- gpio1_s1_translator:av_write -> gpio1_s1_translator_avalon_anti_slave_0_write:in
	signal gpio1_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- gpio1:readdata -> gpio1_s1_translator:av_readdata
	signal vga_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- vga_s1_translator:av_writedata -> vga:avs_s1_writedata
	signal vga_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- vga_s1_translator:av_address -> vga:avs_s1_address
	signal vga_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- vga_s1_translator:av_write -> vga:avs_s1_write
	signal vga_s1_translator_avalon_anti_slave_0_read                                                        : std_logic;                      -- vga_s1_translator:av_read -> vga:avs_s1_read
	signal vga_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- vga:avs_s1_readdata -> vga_s1_translator:av_readdata
	signal blcon_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- blcon_s1_translator:av_writedata -> blcon:writedata
	signal blcon_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- blcon_s1_translator:av_write -> blcon:write
	signal blcon_s1_translator_avalon_anti_slave_0_read                                                      : std_logic;                      -- blcon_s1_translator:av_read -> blcon:read
	signal blcon_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- blcon:readdata -> blcon_s1_translator:av_readdata
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_fast_instruction_master_translator:uav_waitrequest
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(5 downto 0);   -- nios2_fast_instruction_master_translator:uav_burstcount -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0);  -- nios2_fast_instruction_master_translator:uav_writedata -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(31 downto 0);  -- nios2_fast_instruction_master_translator:uav_address -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                      -- nios2_fast_instruction_master_translator:uav_lock -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                      -- nios2_fast_instruction_master_translator:uav_write -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                      -- nios2_fast_instruction_master_translator:uav_read -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0);  -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_fast_instruction_master_translator:uav_readdata
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                      -- nios2_fast_instruction_master_translator:uav_debugaccess -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);   -- nios2_fast_instruction_master_translator:uav_byteenable -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_fast_instruction_master_translator:uav_readdatavalid
	signal nios2_fast_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_fast_data_master_translator:uav_waitrequest
	signal nios2_fast_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(5 downto 0);   -- nios2_fast_data_master_translator:uav_burstcount -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_fast_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_fast_data_master_translator:uav_writedata -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_fast_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(31 downto 0);  -- nios2_fast_data_master_translator:uav_address -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_fast_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                      -- nios2_fast_data_master_translator:uav_lock -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_fast_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                      -- nios2_fast_data_master_translator:uav_write -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_fast_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                      -- nios2_fast_data_master_translator:uav_read -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_fast_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_fast_data_master_translator:uav_readdata
	signal nios2_fast_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                      -- nios2_fast_data_master_translator:uav_debugaccess -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_fast_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_fast_data_master_translator:uav_byteenable -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_fast_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_fast_data_master_translator:uav_readdatavalid
	signal spu_m1_translator_avalon_universal_master_0_waitrequest                                           : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:av_waitrequest -> spu_m1_translator:uav_waitrequest
	signal spu_m1_translator_avalon_universal_master_0_burstcount                                            : std_logic_vector(3 downto 0);   -- spu_m1_translator:uav_burstcount -> spu_m1_translator_avalon_universal_master_0_agent:av_burstcount
	signal spu_m1_translator_avalon_universal_master_0_writedata                                             : std_logic_vector(15 downto 0);  -- spu_m1_translator:uav_writedata -> spu_m1_translator_avalon_universal_master_0_agent:av_writedata
	signal spu_m1_translator_avalon_universal_master_0_address                                               : std_logic_vector(31 downto 0);  -- spu_m1_translator:uav_address -> spu_m1_translator_avalon_universal_master_0_agent:av_address
	signal spu_m1_translator_avalon_universal_master_0_lock                                                  : std_logic;                      -- spu_m1_translator:uav_lock -> spu_m1_translator_avalon_universal_master_0_agent:av_lock
	signal spu_m1_translator_avalon_universal_master_0_write                                                 : std_logic;                      -- spu_m1_translator:uav_write -> spu_m1_translator_avalon_universal_master_0_agent:av_write
	signal spu_m1_translator_avalon_universal_master_0_read                                                  : std_logic;                      -- spu_m1_translator:uav_read -> spu_m1_translator_avalon_universal_master_0_agent:av_read
	signal spu_m1_translator_avalon_universal_master_0_readdata                                              : std_logic_vector(15 downto 0);  -- spu_m1_translator_avalon_universal_master_0_agent:av_readdata -> spu_m1_translator:uav_readdata
	signal spu_m1_translator_avalon_universal_master_0_debugaccess                                           : std_logic;                      -- spu_m1_translator:uav_debugaccess -> spu_m1_translator_avalon_universal_master_0_agent:av_debugaccess
	signal spu_m1_translator_avalon_universal_master_0_byteenable                                            : std_logic_vector(1 downto 0);   -- spu_m1_translator:uav_byteenable -> spu_m1_translator_avalon_universal_master_0_agent:av_byteenable
	signal spu_m1_translator_avalon_universal_master_0_readdatavalid                                         : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:av_readdatavalid -> spu_m1_translator:uav_readdatavalid
	signal vga_m1_translator_avalon_universal_master_0_waitrequest                                           : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:av_waitrequest -> vga_m1_translator:uav_waitrequest
	signal vga_m1_translator_avalon_universal_master_0_burstcount                                            : std_logic_vector(11 downto 0);  -- vga_m1_translator:uav_burstcount -> vga_m1_translator_avalon_universal_master_0_agent:av_burstcount
	signal vga_m1_translator_avalon_universal_master_0_writedata                                             : std_logic_vector(31 downto 0);  -- vga_m1_translator:uav_writedata -> vga_m1_translator_avalon_universal_master_0_agent:av_writedata
	signal vga_m1_translator_avalon_universal_master_0_address                                               : std_logic_vector(31 downto 0);  -- vga_m1_translator:uav_address -> vga_m1_translator_avalon_universal_master_0_agent:av_address
	signal vga_m1_translator_avalon_universal_master_0_lock                                                  : std_logic;                      -- vga_m1_translator:uav_lock -> vga_m1_translator_avalon_universal_master_0_agent:av_lock
	signal vga_m1_translator_avalon_universal_master_0_write                                                 : std_logic;                      -- vga_m1_translator:uav_write -> vga_m1_translator_avalon_universal_master_0_agent:av_write
	signal vga_m1_translator_avalon_universal_master_0_read                                                  : std_logic;                      -- vga_m1_translator:uav_read -> vga_m1_translator_avalon_universal_master_0_agent:av_read
	signal vga_m1_translator_avalon_universal_master_0_readdata                                              : std_logic_vector(31 downto 0);  -- vga_m1_translator_avalon_universal_master_0_agent:av_readdata -> vga_m1_translator:uav_readdata
	signal vga_m1_translator_avalon_universal_master_0_debugaccess                                           : std_logic;                      -- vga_m1_translator:uav_debugaccess -> vga_m1_translator_avalon_universal_master_0_agent:av_debugaccess
	signal vga_m1_translator_avalon_universal_master_0_byteenable                                            : std_logic_vector(3 downto 0);   -- vga_m1_translator:uav_byteenable -> vga_m1_translator_avalon_universal_master_0_agent:av_byteenable
	signal vga_m1_translator_avalon_universal_master_0_readdatavalid                                         : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:av_readdatavalid -> vga_m1_translator:uav_readdatavalid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- nios2_fast_jtag_debug_module_translator:uav_waitrequest -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_fast_jtag_debug_module_translator:uav_burstcount
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_fast_jtag_debug_module_translator:uav_writedata
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0);  -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_fast_jtag_debug_module_translator:uav_address
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_fast_jtag_debug_module_translator:uav_write
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_fast_jtag_debug_module_translator:uav_lock
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_fast_jtag_debug_module_translator:uav_read
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- nios2_fast_jtag_debug_module_translator:uav_readdata -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- nios2_fast_jtag_debug_module_translator:uav_readdatavalid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_fast_jtag_debug_module_translator:uav_debugaccess
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_fast_jtag_debug_module_translator:uav_byteenable
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(115 downto 0); -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(115 downto 0); -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(33 downto 0);  -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                            : std_logic;                      -- ipl_memory_s1_translator:uav_waitrequest -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                             : std_logic_vector(2 downto 0);   -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ipl_memory_s1_translator:uav_burstcount
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                              : std_logic_vector(31 downto 0);  -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ipl_memory_s1_translator:uav_writedata
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                                : std_logic_vector(31 downto 0);  -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> ipl_memory_s1_translator:uav_address
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                                  : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> ipl_memory_s1_translator:uav_write
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                   : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ipl_memory_s1_translator:uav_lock
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                   : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> ipl_memory_s1_translator:uav_read
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                               : std_logic_vector(31 downto 0);  -- ipl_memory_s1_translator:uav_readdata -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                          : std_logic;                      -- ipl_memory_s1_translator:uav_readdatavalid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                            : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ipl_memory_s1_translator:uav_debugaccess
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                             : std_logic_vector(3 downto 0);   -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ipl_memory_s1_translator:uav_byteenable
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                     : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                           : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                   : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                            : std_logic_vector(115 downto 0); -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                           : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                  : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                        : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                         : std_logic_vector(115 downto 0); -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                        : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                      : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                       : std_logic_vector(33 downto 0);  -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                      : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                      : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                       : std_logic_vector(33 downto 0);  -- ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                      : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(15 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(31 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(15 downto 0);  -- sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(97 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(97 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                            : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- peripherals_bridge_s0_translator:uav_waitrequest -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> peripherals_bridge_s0_translator:uav_burstcount
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> peripherals_bridge_s0_translator:uav_writedata
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(31 downto 0);  -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> peripherals_bridge_s0_translator:uav_address
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> peripherals_bridge_s0_translator:uav_write
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> peripherals_bridge_s0_translator:uav_lock
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> peripherals_bridge_s0_translator:uav_read
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- peripherals_bridge_s0_translator:uav_readdata -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- peripherals_bridge_s0_translator:uav_readdatavalid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> peripherals_bridge_s0_translator:uav_debugaccess
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> peripherals_bridge_s0_translator:uav_byteenable
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(115 downto 0); -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(115 downto 0); -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid              : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data               : std_logic_vector(33 downto 0);  -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready              : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> peripherals_bridge_m0_translator:uav_waitrequest
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(2 downto 0);   -- peripherals_bridge_m0_translator:uav_burstcount -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_writedata                              : std_logic_vector(31 downto 0);  -- peripherals_bridge_m0_translator:uav_writedata -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_address                                : std_logic_vector(13 downto 0);  -- peripherals_bridge_m0_translator:uav_address -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- peripherals_bridge_m0_translator:uav_lock -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_write                                  : std_logic;                      -- peripherals_bridge_m0_translator:uav_write -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_read                                   : std_logic;                      -- peripherals_bridge_m0_translator:uav_read -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_readdata                               : std_logic_vector(31 downto 0);  -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> peripherals_bridge_m0_translator:uav_readdata
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- peripherals_bridge_m0_translator:uav_debugaccess -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(3 downto 0);   -- peripherals_bridge_m0_translator:uav_byteenable -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> peripherals_bridge_m0_translator:uav_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(13 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(87 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(87 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                      -- sysuart_s1_translator:uav_waitrequest -> sysuart_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);   -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysuart_s1_translator:uav_burstcount
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sysuart_s1_translator:uav_writedata
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(13 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_address -> sysuart_s1_translator:uav_address
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_write -> sysuart_s1_translator:uav_write
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sysuart_s1_translator:uav_lock
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_read -> sysuart_s1_translator:uav_read
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0);  -- sysuart_s1_translator:uav_readdata -> sysuart_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                      -- sysuart_s1_translator:uav_readdatavalid -> sysuart_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysuart_s1_translator:uav_debugaccess
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);   -- sysuart_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysuart_s1_translator:uav_byteenable
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(87 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysuart_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysuart_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(87 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysuart_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysuart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(13 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(87 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(87 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                      -- systimer_s1_translator:uav_waitrequest -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);   -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> systimer_s1_translator:uav_burstcount
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> systimer_s1_translator:uav_writedata
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(13 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_address -> systimer_s1_translator:uav_address
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_write -> systimer_s1_translator:uav_write
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> systimer_s1_translator:uav_lock
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_read -> systimer_s1_translator:uav_read
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0);  -- systimer_s1_translator:uav_readdata -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                      -- systimer_s1_translator:uav_readdatavalid -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> systimer_s1_translator:uav_debugaccess
	signal systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);   -- systimer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> systimer_s1_translator:uav_byteenable
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(87 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(87 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(33 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(13 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(87 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(87 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                      -- led_7seg_s1_translator:uav_waitrequest -> led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);   -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_7seg_s1_translator:uav_burstcount
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_7seg_s1_translator:uav_writedata
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(13 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_7seg_s1_translator:uav_address
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_7seg_s1_translator:uav_write
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_7seg_s1_translator:uav_lock
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_7seg_s1_translator:uav_read
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0);  -- led_7seg_s1_translator:uav_readdata -> led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                      -- led_7seg_s1_translator:uav_readdatavalid -> led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_7seg_s1_translator:uav_debugaccess
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);   -- led_7seg_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_7seg_s1_translator:uav_byteenable
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(87 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(87 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(33 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- psw_s1_translator:uav_waitrequest -> psw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- psw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> psw_s1_translator:uav_burstcount
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> psw_s1_translator:uav_writedata
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(13 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent:m0_address -> psw_s1_translator:uav_address
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:m0_write -> psw_s1_translator:uav_write
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> psw_s1_translator:uav_lock
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:m0_read -> psw_s1_translator:uav_read
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- psw_s1_translator:uav_readdata -> psw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- psw_s1_translator:uav_readdatavalid -> psw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> psw_s1_translator:uav_debugaccess
	signal psw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- psw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> psw_s1_translator:uav_byteenable
	signal psw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal psw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(87 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal psw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> psw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> psw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> psw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> psw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(87 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> psw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> psw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- dipsw_s1_translator:uav_waitrequest -> dipsw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dipsw_s1_translator:uav_burstcount
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dipsw_s1_translator:uav_writedata
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(13 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_address -> dipsw_s1_translator:uav_address
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_write -> dipsw_s1_translator:uav_write
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dipsw_s1_translator:uav_lock
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_read -> dipsw_s1_translator:uav_read
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- dipsw_s1_translator:uav_readdata -> dipsw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- dipsw_s1_translator:uav_readdatavalid -> dipsw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dipsw_s1_translator:uav_debugaccess
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- dipsw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dipsw_s1_translator:uav_byteenable
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(87 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dipsw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dipsw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(87 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dipsw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dipsw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- spu_s1_translator:uav_waitrequest -> spu_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- spu_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> spu_s1_translator:uav_burstcount
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> spu_s1_translator:uav_writedata
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(13 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent:m0_address -> spu_s1_translator:uav_address
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:m0_write -> spu_s1_translator:uav_write
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:m0_lock -> spu_s1_translator:uav_lock
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:m0_read -> spu_s1_translator:uav_read
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- spu_s1_translator:uav_readdata -> spu_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- spu_s1_translator:uav_readdatavalid -> spu_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spu_s1_translator:uav_debugaccess
	signal spu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- spu_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> spu_s1_translator:uav_byteenable
	signal spu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal spu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(87 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal spu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spu_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spu_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spu_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spu_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(87 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spu_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spu_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                      -- mmcdma_s1_translator:uav_waitrequest -> mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);   -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mmcdma_s1_translator:uav_burstcount
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mmcdma_s1_translator:uav_writedata
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(13 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_address -> mmcdma_s1_translator:uav_address
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_write -> mmcdma_s1_translator:uav_write
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mmcdma_s1_translator:uav_lock
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_read -> mmcdma_s1_translator:uav_read
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0);  -- mmcdma_s1_translator:uav_readdata -> mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                      -- mmcdma_s1_translator:uav_readdatavalid -> mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mmcdma_s1_translator:uav_debugaccess
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);   -- mmcdma_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mmcdma_s1_translator:uav_byteenable
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(87 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(87 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- ps2_keyboard_avalon_slave_translator:uav_waitrequest -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ps2_keyboard_avalon_slave_translator:uav_burstcount
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ps2_keyboard_avalon_slave_translator:uav_writedata
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(13 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> ps2_keyboard_avalon_slave_translator:uav_address
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> ps2_keyboard_avalon_slave_translator:uav_write
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ps2_keyboard_avalon_slave_translator:uav_lock
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> ps2_keyboard_avalon_slave_translator:uav_read
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- ps2_keyboard_avalon_slave_translator:uav_readdata -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- ps2_keyboard_avalon_slave_translator:uav_readdatavalid -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ps2_keyboard_avalon_slave_translator:uav_debugaccess
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ps2_keyboard_avalon_slave_translator:uav_byteenable
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(87 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(87 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- gpio1_s1_translator:uav_waitrequest -> gpio1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> gpio1_s1_translator:uav_burstcount
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> gpio1_s1_translator:uav_writedata
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(13 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_address -> gpio1_s1_translator:uav_address
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_write -> gpio1_s1_translator:uav_write
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> gpio1_s1_translator:uav_lock
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_read -> gpio1_s1_translator:uav_read
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- gpio1_s1_translator:uav_readdata -> gpio1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- gpio1_s1_translator:uav_readdatavalid -> gpio1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gpio1_s1_translator:uav_debugaccess
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- gpio1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> gpio1_s1_translator:uav_byteenable
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(87 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gpio1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gpio1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(87 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gpio1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gpio1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- vga_s1_translator:uav_waitrequest -> vga_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- vga_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> vga_s1_translator:uav_burstcount
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> vga_s1_translator:uav_writedata
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(13 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent:m0_address -> vga_s1_translator:uav_address
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:m0_write -> vga_s1_translator:uav_write
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:m0_lock -> vga_s1_translator:uav_lock
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:m0_read -> vga_s1_translator:uav_read
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- vga_s1_translator:uav_readdata -> vga_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- vga_s1_translator:uav_readdatavalid -> vga_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> vga_s1_translator:uav_debugaccess
	signal vga_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- vga_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> vga_s1_translator:uav_byteenable
	signal vga_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal vga_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(87 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal vga_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> vga_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> vga_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> vga_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> vga_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(87 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> vga_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> vga_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- blcon_s1_translator:uav_waitrequest -> blcon_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> blcon_s1_translator:uav_burstcount
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> blcon_s1_translator:uav_writedata
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(13 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_address -> blcon_s1_translator:uav_address
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_write -> blcon_s1_translator:uav_write
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_lock -> blcon_s1_translator:uav_lock
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_read -> blcon_s1_translator:uav_read
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- blcon_s1_translator:uav_readdata -> blcon_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- blcon_s1_translator:uav_readdatavalid -> blcon_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> blcon_s1_translator:uav_debugaccess
	signal blcon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- blcon_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> blcon_s1_translator:uav_byteenable
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(87 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> blcon_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> blcon_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(87 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> blcon_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> blcon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(114 downto 0); -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                      -- addr_router:sink_ready -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(114 downto 0); -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                      -- addr_router_001:sink_ready -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal spu_m1_translator_avalon_universal_master_0_agent_cp_endofpacket                                  : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal spu_m1_translator_avalon_universal_master_0_agent_cp_valid                                        : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal spu_m1_translator_avalon_universal_master_0_agent_cp_startofpacket                                : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal spu_m1_translator_avalon_universal_master_0_agent_cp_data                                         : std_logic_vector(96 downto 0);  -- spu_m1_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal spu_m1_translator_avalon_universal_master_0_agent_cp_ready                                        : std_logic;                      -- addr_router_002:sink_ready -> spu_m1_translator_avalon_universal_master_0_agent:cp_ready
	signal vga_m1_translator_avalon_universal_master_0_agent_cp_endofpacket                                  : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	signal vga_m1_translator_avalon_universal_master_0_agent_cp_valid                                        : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	signal vga_m1_translator_avalon_universal_master_0_agent_cp_startofpacket                                : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	signal vga_m1_translator_avalon_universal_master_0_agent_cp_data                                         : std_logic_vector(114 downto 0); -- vga_m1_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	signal vga_m1_translator_avalon_universal_master_0_agent_cp_ready                                        : std_logic;                      -- addr_router_003:sink_ready -> vga_m1_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(114 downto 0); -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router:sink_ready -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                            : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                                  : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                          : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                   : std_logic_vector(114 downto 0); -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                                  : std_logic;                      -- id_router_001:sink_ready -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(96 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(114 downto 0); -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_003:sink_ready -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(86 downto 0);  -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	signal peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router_004:sink_ready -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(86 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                      -- id_router_004:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(86 downto 0);  -- sysuart_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal sysuart_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                      -- id_router_005:sink_ready -> sysuart_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(86 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_006:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(86 downto 0);  -- systimer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                      -- id_router_007:sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(86 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_008:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(86 downto 0);  -- led_7seg_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                      -- id_router_009:sink_ready -> led_7seg_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal psw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal psw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal psw_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(86 downto 0);  -- psw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal psw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_010:sink_ready -> psw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(86 downto 0);  -- dipsw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal dipsw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_011:sink_ready -> dipsw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal spu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal spu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal spu_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(86 downto 0);  -- spu_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal spu_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_012:sink_ready -> spu_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(86 downto 0);  -- mmcdma_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                      -- id_router_013:sink_ready -> mmcdma_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(86 downto 0);  -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_014:sink_ready -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(86 downto 0);  -- gpio1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal gpio1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_015:sink_ready -> gpio1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal vga_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal vga_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal vga_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(86 downto 0);  -- vga_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal vga_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_016:sink_ready -> vga_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(86 downto 0);  -- blcon_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	signal blcon_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_017:sink_ready -> blcon_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                       : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                             : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                     : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                              : std_logic_vector(114 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                             : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                       : std_logic;                      -- limiter:rsp_src_endofpacket -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                             : std_logic;                      -- limiter:rsp_src_valid -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                     : std_logic;                      -- limiter:rsp_src_startofpacket -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                              : std_logic_vector(114 downto 0); -- limiter:rsp_src_data -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                           : std_logic_vector(3 downto 0);   -- limiter:rsp_src_channel -> nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                             : std_logic;                      -- nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                                   : std_logic;                      -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                         : std_logic;                      -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                 : std_logic;                      -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                          : std_logic_vector(114 downto 0); -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                       : std_logic_vector(3 downto 0);   -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                         : std_logic;                      -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                                   : std_logic;                      -- limiter_001:rsp_src_endofpacket -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                         : std_logic;                      -- limiter_001:rsp_src_valid -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_001_rsp_src_startofpacket                                                                 : std_logic;                      -- limiter_001:rsp_src_startofpacket -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_001_rsp_src_data                                                                          : std_logic_vector(114 downto 0); -- limiter_001:rsp_src_data -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_001_rsp_src_channel                                                                       : std_logic_vector(3 downto 0);   -- limiter_001:rsp_src_channel -> nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_001_rsp_src_ready                                                                         : std_logic;                      -- nios2_fast_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	signal addr_router_004_src_endofpacket                                                                   : std_logic;                      -- addr_router_004:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	signal addr_router_004_src_valid                                                                         : std_logic;                      -- addr_router_004:src_valid -> limiter_002:cmd_sink_valid
	signal addr_router_004_src_startofpacket                                                                 : std_logic;                      -- addr_router_004:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	signal addr_router_004_src_data                                                                          : std_logic_vector(86 downto 0);  -- addr_router_004:src_data -> limiter_002:cmd_sink_data
	signal addr_router_004_src_channel                                                                       : std_logic_vector(13 downto 0);  -- addr_router_004:src_channel -> limiter_002:cmd_sink_channel
	signal addr_router_004_src_ready                                                                         : std_logic;                      -- limiter_002:cmd_sink_ready -> addr_router_004:src_ready
	signal limiter_002_rsp_src_endofpacket                                                                   : std_logic;                      -- limiter_002:rsp_src_endofpacket -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_002_rsp_src_valid                                                                         : std_logic;                      -- limiter_002:rsp_src_valid -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_002_rsp_src_startofpacket                                                                 : std_logic;                      -- limiter_002:rsp_src_startofpacket -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_002_rsp_src_data                                                                          : std_logic_vector(86 downto 0);  -- limiter_002:rsp_src_data -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_002_rsp_src_channel                                                                       : std_logic_vector(13 downto 0);  -- limiter_002:rsp_src_channel -> peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_002_rsp_src_ready                                                                         : std_logic;                      -- peripherals_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                 : std_logic;                      -- burst_adapter:source0_endofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                       : std_logic;                      -- burst_adapter:source0_valid -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                               : std_logic;                      -- burst_adapter:source0_startofpacket -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                        : std_logic_vector(114 downto 0); -- burst_adapter:source0_data -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                       : std_logic;                      -- nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                     : std_logic_vector(3 downto 0);   -- burst_adapter:source0_channel -> nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                             : std_logic;                      -- burst_adapter_001:source0_endofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                   : std_logic;                      -- burst_adapter_001:source0_valid -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                           : std_logic;                      -- burst_adapter_001:source0_startofpacket -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                    : std_logic_vector(114 downto 0); -- burst_adapter_001:source0_data -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                   : std_logic;                      -- ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                 : std_logic_vector(3 downto 0);   -- burst_adapter_001:source0_channel -> ipl_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_002_source0_endofpacket                                                             : std_logic;                      -- burst_adapter_002:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_002_source0_valid                                                                   : std_logic;                      -- burst_adapter_002:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_002_source0_startofpacket                                                           : std_logic;                      -- burst_adapter_002:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_002_source0_data                                                                    : std_logic_vector(96 downto 0);  -- burst_adapter_002:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_002_source0_ready                                                                   : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	signal burst_adapter_002_source0_channel                                                                 : std_logic_vector(3 downto 0);   -- burst_adapter_002:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_003_source0_endofpacket                                                             : std_logic;                      -- burst_adapter_003:source0_endofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_003_source0_valid                                                                   : std_logic;                      -- burst_adapter_003:source0_valid -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_003_source0_startofpacket                                                           : std_logic;                      -- burst_adapter_003:source0_startofpacket -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_003_source0_data                                                                    : std_logic_vector(114 downto 0); -- burst_adapter_003:source0_data -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_003_source0_ready                                                                   : std_logic;                      -- peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	signal burst_adapter_003_source0_channel                                                                 : std_logic_vector(3 downto 0);   -- burst_adapter_003:source0_channel -> peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                    : std_logic;                      -- rst_controller:reset_out -> [addr_router_004:reset, blcon:reset, blcon_s1_translator:reset, blcon_s1_translator_avalon_universal_slave_0_agent:reset, blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_004:reset, dipsw_s1_translator:reset, dipsw_s1_translator_avalon_universal_slave_0_agent:reset, dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, gpio1_s1_translator:reset, gpio1_s1_translator_avalon_universal_slave_0_agent:reset, gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_7seg_s1_translator:reset, led_7seg_s1_translator_avalon_universal_slave_0_agent:reset, led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, mmcdma:reset, mmcdma_s1_translator:reset, mmcdma_s1_translator_avalon_universal_slave_0_agent:reset, mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, peripherals_bridge:m0_reset, peripherals_bridge_m0_translator:reset, peripherals_bridge_m0_translator_avalon_universal_master_0_agent:reset, ps2_keyboard:reset, ps2_keyboard_avalon_slave_translator:reset, ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:reset, ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, psw_s1_translator:reset, psw_s1_translator_avalon_universal_slave_0_agent:reset, psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_mux_004:reset, rst_controller_reset_out_reset:in, spu:csi_global_reset, spu_s1_translator:reset, spu_s1_translator_avalon_universal_slave_0_agent:reset, spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, systimer_s1_translator:reset, systimer_s1_translator_avalon_universal_slave_0_agent:reset, systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysuart_s1_translator:reset, sysuart_s1_translator_avalon_universal_slave_0_agent:reset, sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, vga:g_reset, vga_s1_translator:reset, vga_s1_translator_avalon_universal_slave_0_agent:reset, vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal rst_controller_001_reset_out_reset                                                                : std_logic;                      -- rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, ipl_memory:reset, ipl_memory_s1_translator:reset, ipl_memory_s1_translator_avalon_universal_slave_0_agent:reset, ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, limiter:reset, limiter_001:reset, nios2_fast_data_master_translator:reset, nios2_fast_data_master_translator_avalon_universal_master_0_agent:reset, nios2_fast_instruction_master_translator:reset, nios2_fast_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_fast_jtag_debug_module_translator:reset, nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, peripherals_bridge:s0_reset, peripherals_bridge_s0_translator:reset, peripherals_bridge_s0_translator_avalon_universal_slave_0_agent:reset, peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_001_reset_out_reset:in, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	signal rst_controller_001_reset_out_reset_req                                                            : std_logic;                      -- rst_controller_001:reset_req -> ipl_memory:reset_req
	signal rst_controller_002_reset_out_reset                                                                : std_logic;                      -- rst_controller_002:reset_out -> [addr_router_002:reset, addr_router_003:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, spu_m1_translator:reset, spu_m1_translator_avalon_universal_master_0_agent:reset, vga_m1_translator:reset, vga_m1_translator_avalon_universal_master_0_agent:reset, width_adapter_002:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                          : std_logic_vector(114 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                         : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                          : std_logic_vector(114 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                         : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                     : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                      : std_logic_vector(114 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                     : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                     : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                      : std_logic_vector(114 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                     : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> burst_adapter_003:sink0_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                     : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> burst_adapter_003:sink0_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> burst_adapter_003:sink0_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                      : std_logic_vector(114 downto 0); -- cmd_xbar_demux_001:src3_data -> burst_adapter_003:sink0_data
	signal cmd_xbar_demux_001_src3_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src3_channel -> burst_adapter_003:sink0_channel
	signal cmd_xbar_demux_002_src0_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                     : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_002:sink2_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                      : std_logic_vector(96 downto 0);  -- cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_002:sink2_data
	signal cmd_xbar_demux_002_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_002:sink2_channel
	signal cmd_xbar_demux_002_src0_ready                                                                     : std_logic;                      -- cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                          : std_logic_vector(114 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                          : std_logic_vector(114 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                         : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                      : std_logic_vector(114 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                     : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                      : std_logic_vector(114 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                     : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src2_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src2_endofpacket -> spu_m1_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_002_src2_valid                                                                     : std_logic;                      -- rsp_xbar_demux_002:src2_valid -> spu_m1_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_002_src2_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_002:src2_startofpacket -> spu_m1_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_002_src2_data                                                                      : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_002:src2_data -> spu_m1_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_002_src2_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_002:src2_channel -> spu_m1_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_003_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                      : std_logic_vector(114 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal limiter_cmd_src_endofpacket                                                                       : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                     : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                              : std_logic_vector(114 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                           : std_logic_vector(3 downto 0);   -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                      : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                            : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                    : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                             : std_logic_vector(114 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                          : std_logic_vector(3 downto 0);   -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                            : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                                   : std_logic;                      -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                                 : std_logic;                      -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                          : std_logic_vector(114 downto 0); -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                       : std_logic_vector(3 downto 0);   -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                         : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                  : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                        : std_logic;                      -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                         : std_logic_vector(114 downto 0); -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                      : std_logic_vector(3 downto 0);   -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                        : std_logic;                      -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal addr_router_002_src_endofpacket                                                                   : std_logic;                      -- addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal addr_router_002_src_valid                                                                         : std_logic;                      -- addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	signal addr_router_002_src_startofpacket                                                                 : std_logic;                      -- addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal addr_router_002_src_data                                                                          : std_logic_vector(96 downto 0);  -- addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	signal addr_router_002_src_channel                                                                       : std_logic_vector(3 downto 0);   -- addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	signal addr_router_002_src_ready                                                                         : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	signal rsp_xbar_demux_002_src2_ready                                                                     : std_logic;                      -- spu_m1_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_002:src2_ready
	signal addr_router_003_src_endofpacket                                                                   : std_logic;                      -- addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	signal addr_router_003_src_valid                                                                         : std_logic;                      -- addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	signal addr_router_003_src_startofpacket                                                                 : std_logic;                      -- addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	signal addr_router_003_src_data                                                                          : std_logic_vector(114 downto 0); -- addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	signal addr_router_003_src_channel                                                                       : std_logic_vector(3 downto 0);   -- addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	signal addr_router_003_src_ready                                                                         : std_logic;                      -- cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	signal width_adapter_005_src_ready                                                                       : std_logic;                      -- vga_m1_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_005:out_ready
	signal cmd_xbar_mux_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_src_data                                                                             : std_logic_vector(114 downto 0); -- cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_src_channel                                                                          : std_logic_vector(3 downto 0);   -- cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_src_ready                                                                            : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                         : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                               : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                       : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                : std_logic_vector(114 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                             : std_logic_vector(3 downto 0);   -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                        : std_logic;                      -- cmd_xbar_mux_001:src_valid -> burst_adapter_001:sink0_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                         : std_logic_vector(114 downto 0); -- cmd_xbar_mux_001:src_data -> burst_adapter_001:sink0_data
	signal cmd_xbar_mux_001_src_channel                                                                      : std_logic_vector(3 downto 0);   -- cmd_xbar_mux_001:src_channel -> burst_adapter_001:sink0_channel
	signal cmd_xbar_mux_001_src_ready                                                                        : std_logic;                      -- burst_adapter_001:sink0_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                     : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                           : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                   : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                            : std_logic_vector(114 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                         : std_logic_vector(3 downto 0);   -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                        : std_logic;                      -- cmd_xbar_mux_002:src_valid -> burst_adapter_002:sink0_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                         : std_logic_vector(96 downto 0);  -- cmd_xbar_mux_002:src_data -> burst_adapter_002:sink0_data
	signal cmd_xbar_mux_002_src_channel                                                                      : std_logic_vector(3 downto 0);   -- cmd_xbar_mux_002:src_channel -> burst_adapter_002:sink0_channel
	signal cmd_xbar_mux_002_src_ready                                                                        : std_logic;                      -- burst_adapter_002:sink0_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                     : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                           : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                   : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                            : std_logic_vector(96 downto 0);  -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                         : std_logic_vector(3 downto 0);   -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_001_src3_ready                                                                     : std_logic;                      -- burst_adapter_003:sink0_ready -> cmd_xbar_demux_001:src3_ready
	signal id_router_003_src_endofpacket                                                                     : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                           : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                   : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                            : std_logic_vector(114 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                         : std_logic_vector(3 downto 0);   -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_004_src0_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src0_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src0_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src0_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src1_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src1_endofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src1_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src1_valid -> sysuart_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src1_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src1_startofpacket -> sysuart_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src1_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src1_data -> sysuart_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src1_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src1_channel -> sysuart_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src2_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src2_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src2_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src2_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src2_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src2_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src2_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src2_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src2_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src2_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src3_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src3_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src3_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src3_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src3_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src3_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src3_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src3_data -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src3_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src3_channel -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src4_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src4_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src4_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src4_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src4_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src4_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src4_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src4_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src4_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src4_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src5_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src5_endofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src5_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src5_valid -> led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src5_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src5_startofpacket -> led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src5_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src5_data -> led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src5_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src5_channel -> led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src6_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src6_endofpacket -> psw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src6_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src6_valid -> psw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src6_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src6_startofpacket -> psw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src6_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src6_data -> psw_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src6_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src6_channel -> psw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src7_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src7_endofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src7_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src7_valid -> dipsw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src7_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src7_startofpacket -> dipsw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src7_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src7_data -> dipsw_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src7_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src7_channel -> dipsw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src8_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src8_endofpacket -> spu_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src8_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src8_valid -> spu_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src8_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src8_startofpacket -> spu_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src8_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src8_data -> spu_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src8_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src8_channel -> spu_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src9_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_004:src9_endofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src9_valid                                                                     : std_logic;                      -- cmd_xbar_demux_004:src9_valid -> mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src9_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_004:src9_startofpacket -> mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src9_data                                                                      : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src9_data -> mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src9_channel                                                                   : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src9_channel -> mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src10_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux_004:src10_endofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src10_valid                                                                    : std_logic;                      -- cmd_xbar_demux_004:src10_valid -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src10_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux_004:src10_startofpacket -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src10_data                                                                     : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src10_data -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src10_channel                                                                  : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src10_channel -> ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src11_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux_004:src11_endofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src11_valid                                                                    : std_logic;                      -- cmd_xbar_demux_004:src11_valid -> gpio1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src11_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux_004:src11_startofpacket -> gpio1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src11_data                                                                     : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src11_data -> gpio1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src11_channel                                                                  : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src11_channel -> gpio1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src12_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux_004:src12_endofpacket -> vga_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src12_valid                                                                    : std_logic;                      -- cmd_xbar_demux_004:src12_valid -> vga_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src12_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux_004:src12_startofpacket -> vga_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src12_data                                                                     : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src12_data -> vga_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src12_channel                                                                  : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src12_channel -> vga_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_004_src13_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux_004:src13_endofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_004_src13_valid                                                                    : std_logic;                      -- cmd_xbar_demux_004:src13_valid -> blcon_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_004_src13_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux_004:src13_startofpacket -> blcon_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_004_src13_data                                                                     : std_logic_vector(86 downto 0);  -- cmd_xbar_demux_004:src13_data -> blcon_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_004_src13_channel                                                                  : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_004:src13_channel -> blcon_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_004_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_004:sink0_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_004:sink0_data
	signal rsp_xbar_demux_004_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_004:sink0_channel
	signal rsp_xbar_demux_004_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_004:sink1_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_004:sink1_data
	signal rsp_xbar_demux_005_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_004:sink1_channel
	signal rsp_xbar_demux_005_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink1_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_004:sink2_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_004:sink2_data
	signal rsp_xbar_demux_006_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_004:sink2_channel
	signal rsp_xbar_demux_006_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_004:sink3_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_004:sink3_data
	signal rsp_xbar_demux_007_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_004:sink3_channel
	signal rsp_xbar_demux_007_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink3_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_004:sink4_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_004:sink4_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_004:sink4_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_004:sink4_data
	signal rsp_xbar_demux_008_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_004:sink4_channel
	signal rsp_xbar_demux_008_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink4_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_004:sink5_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_004:sink5_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_004:sink5_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_004:sink5_data
	signal rsp_xbar_demux_009_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_004:sink5_channel
	signal rsp_xbar_demux_009_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink5_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_004:sink6_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_004:sink6_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_004:sink6_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_004:sink6_data
	signal rsp_xbar_demux_010_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_004:sink6_channel
	signal rsp_xbar_demux_010_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink6_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_004:sink7_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_004:sink7_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_004:sink7_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_004:sink7_data
	signal rsp_xbar_demux_011_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_004:sink7_channel
	signal rsp_xbar_demux_011_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink7_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_004:sink8_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_004:sink8_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_004:sink8_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_004:sink8_data
	signal rsp_xbar_demux_012_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_004:sink8_channel
	signal rsp_xbar_demux_012_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink8_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_004:sink9_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_004:sink9_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_004:sink9_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_004:sink9_data
	signal rsp_xbar_demux_013_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_004:sink9_channel
	signal rsp_xbar_demux_013_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink9_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_004:sink10_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_004:sink10_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_004:sink10_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_004:sink10_data
	signal rsp_xbar_demux_014_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_004:sink10_channel
	signal rsp_xbar_demux_014_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink10_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_004:sink11_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_004:sink11_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_004:sink11_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_004:sink11_data
	signal rsp_xbar_demux_015_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_004:sink11_channel
	signal rsp_xbar_demux_015_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink11_ready -> rsp_xbar_demux_015:src0_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_004:sink12_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_004:sink12_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_004:sink12_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_004:sink12_data
	signal rsp_xbar_demux_016_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_004:sink12_channel
	signal rsp_xbar_demux_016_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink12_ready -> rsp_xbar_demux_016:src0_ready
	signal rsp_xbar_demux_017_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_004:sink13_endofpacket
	signal rsp_xbar_demux_017_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_004:sink13_valid
	signal rsp_xbar_demux_017_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_004:sink13_startofpacket
	signal rsp_xbar_demux_017_src0_data                                                                      : std_logic_vector(86 downto 0);  -- rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_004:sink13_data
	signal rsp_xbar_demux_017_src0_channel                                                                   : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_004:sink13_channel
	signal rsp_xbar_demux_017_src0_ready                                                                     : std_logic;                      -- rsp_xbar_mux_004:sink13_ready -> rsp_xbar_demux_017:src0_ready
	signal limiter_002_cmd_src_endofpacket                                                                   : std_logic;                      -- limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	signal limiter_002_cmd_src_startofpacket                                                                 : std_logic;                      -- limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	signal limiter_002_cmd_src_data                                                                          : std_logic_vector(86 downto 0);  -- limiter_002:cmd_src_data -> cmd_xbar_demux_004:sink_data
	signal limiter_002_cmd_src_channel                                                                       : std_logic_vector(13 downto 0);  -- limiter_002:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	signal limiter_002_cmd_src_ready                                                                         : std_logic;                      -- cmd_xbar_demux_004:sink_ready -> limiter_002:cmd_src_ready
	signal rsp_xbar_mux_004_src_endofpacket                                                                  : std_logic;                      -- rsp_xbar_mux_004:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	signal rsp_xbar_mux_004_src_valid                                                                        : std_logic;                      -- rsp_xbar_mux_004:src_valid -> limiter_002:rsp_sink_valid
	signal rsp_xbar_mux_004_src_startofpacket                                                                : std_logic;                      -- rsp_xbar_mux_004:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	signal rsp_xbar_mux_004_src_data                                                                         : std_logic_vector(86 downto 0);  -- rsp_xbar_mux_004:src_data -> limiter_002:rsp_sink_data
	signal rsp_xbar_mux_004_src_channel                                                                      : std_logic_vector(13 downto 0);  -- rsp_xbar_mux_004:src_channel -> limiter_002:rsp_sink_channel
	signal rsp_xbar_mux_004_src_ready                                                                        : std_logic;                      -- limiter_002:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	signal cmd_xbar_demux_004_src0_ready                                                                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src0_ready
	signal id_router_004_src_endofpacket                                                                     : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                           : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                   : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_004_src1_ready                                                                     : std_logic;                      -- sysuart_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src1_ready
	signal id_router_005_src_endofpacket                                                                     : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                           : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                   : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_004_src2_ready                                                                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src2_ready
	signal id_router_006_src_endofpacket                                                                     : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                           : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                   : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_004_src3_ready                                                                     : std_logic;                      -- systimer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src3_ready
	signal id_router_007_src_endofpacket                                                                     : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                           : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                   : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_004_src4_ready                                                                     : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src4_ready
	signal id_router_008_src_endofpacket                                                                     : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                           : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                   : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_004_src5_ready                                                                     : std_logic;                      -- led_7seg_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src5_ready
	signal id_router_009_src_endofpacket                                                                     : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                           : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                   : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_004_src6_ready                                                                     : std_logic;                      -- psw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src6_ready
	signal id_router_010_src_endofpacket                                                                     : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                           : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                   : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_004_src7_ready                                                                     : std_logic;                      -- dipsw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src7_ready
	signal id_router_011_src_endofpacket                                                                     : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                           : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                   : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_004_src8_ready                                                                     : std_logic;                      -- spu_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src8_ready
	signal id_router_012_src_endofpacket                                                                     : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                           : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                   : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_004_src9_ready                                                                     : std_logic;                      -- mmcdma_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src9_ready
	signal id_router_013_src_endofpacket                                                                     : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                           : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                   : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_demux_004_src10_ready                                                                    : std_logic;                      -- ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src10_ready
	signal id_router_014_src_endofpacket                                                                     : std_logic;                      -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                           : std_logic;                      -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                                   : std_logic;                      -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_demux_004_src11_ready                                                                    : std_logic;                      -- gpio1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src11_ready
	signal id_router_015_src_endofpacket                                                                     : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                           : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                   : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_demux_004_src12_ready                                                                    : std_logic;                      -- vga_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src12_ready
	signal id_router_016_src_endofpacket                                                                     : std_logic;                      -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                           : std_logic;                      -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                                   : std_logic;                      -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_demux_004_src13_ready                                                                    : std_logic;                      -- blcon_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_004:src13_ready
	signal id_router_017_src_endofpacket                                                                     : std_logic;                      -- id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	signal id_router_017_src_valid                                                                           : std_logic;                      -- id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	signal id_router_017_src_startofpacket                                                                   : std_logic;                      -- id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	signal id_router_017_src_data                                                                            : std_logic_vector(86 downto 0);  -- id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	signal id_router_017_src_channel                                                                         : std_logic_vector(13 downto 0);  -- id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	signal id_router_017_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                         : std_logic;                      -- cmd_xbar_demux:src2_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src2_data                                                                          : std_logic_vector(114 downto 0); -- cmd_xbar_demux:src2_data -> width_adapter:in_data
	signal cmd_xbar_demux_src2_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src2_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_src2_ready                                                                         : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux:src2_ready
	signal width_adapter_src_endofpacket                                                                     : std_logic;                      -- width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal width_adapter_src_valid                                                                           : std_logic;                      -- width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	signal width_adapter_src_startofpacket                                                                   : std_logic;                      -- width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal width_adapter_src_data                                                                            : std_logic_vector(96 downto 0);  -- width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	signal width_adapter_src_ready                                                                           : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                         : std_logic_vector(3 downto 0);   -- width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_001_src2_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> width_adapter_001:in_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                     : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> width_adapter_001:in_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> width_adapter_001:in_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                      : std_logic_vector(114 downto 0); -- cmd_xbar_demux_001:src2_data -> width_adapter_001:in_data
	signal cmd_xbar_demux_001_src2_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src2_channel -> width_adapter_001:in_channel
	signal cmd_xbar_demux_001_src2_ready                                                                     : std_logic;                      -- width_adapter_001:in_ready -> cmd_xbar_demux_001:src2_ready
	signal width_adapter_001_src_endofpacket                                                                 : std_logic;                      -- width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal width_adapter_001_src_valid                                                                       : std_logic;                      -- width_adapter_001:out_valid -> cmd_xbar_mux_002:sink1_valid
	signal width_adapter_001_src_startofpacket                                                               : std_logic;                      -- width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal width_adapter_001_src_data                                                                        : std_logic_vector(96 downto 0);  -- width_adapter_001:out_data -> cmd_xbar_mux_002:sink1_data
	signal width_adapter_001_src_ready                                                                       : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                     : std_logic_vector(3 downto 0);   -- width_adapter_001:out_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_003_src0_endofpacket                                                               : std_logic;                      -- cmd_xbar_demux_003:src0_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_003_src0_valid                                                                     : std_logic;                      -- cmd_xbar_demux_003:src0_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_003_src0_startofpacket                                                             : std_logic;                      -- cmd_xbar_demux_003:src0_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_003_src0_data                                                                      : std_logic_vector(114 downto 0); -- cmd_xbar_demux_003:src0_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_003_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_003:src0_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_003_src0_ready                                                                     : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_demux_003:src0_ready
	signal width_adapter_002_src_endofpacket                                                                 : std_logic;                      -- width_adapter_002:out_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	signal width_adapter_002_src_valid                                                                       : std_logic;                      -- width_adapter_002:out_valid -> cmd_xbar_mux_002:sink3_valid
	signal width_adapter_002_src_startofpacket                                                               : std_logic;                      -- width_adapter_002:out_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	signal width_adapter_002_src_data                                                                        : std_logic_vector(96 downto 0);  -- width_adapter_002:out_data -> cmd_xbar_mux_002:sink3_data
	signal width_adapter_002_src_ready                                                                       : std_logic;                      -- cmd_xbar_mux_002:sink3_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                     : std_logic_vector(3 downto 0);   -- width_adapter_002:out_channel -> cmd_xbar_mux_002:sink3_channel
	signal rsp_xbar_demux_002_src0_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> width_adapter_003:in_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                     : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> width_adapter_003:in_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> width_adapter_003:in_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                      : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_002:src0_data -> width_adapter_003:in_data
	signal rsp_xbar_demux_002_src0_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_002:src0_channel -> width_adapter_003:in_channel
	signal rsp_xbar_demux_002_src0_ready                                                                     : std_logic;                      -- width_adapter_003:in_ready -> rsp_xbar_demux_002:src0_ready
	signal width_adapter_003_src_endofpacket                                                                 : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal width_adapter_003_src_valid                                                                       : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_mux:sink2_valid
	signal width_adapter_003_src_startofpacket                                                               : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal width_adapter_003_src_data                                                                        : std_logic_vector(114 downto 0); -- width_adapter_003:out_data -> rsp_xbar_mux:sink2_data
	signal width_adapter_003_src_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink2_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                     : std_logic_vector(3 downto 0);   -- width_adapter_003:out_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src1_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> width_adapter_004:in_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                     : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> width_adapter_004:in_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> width_adapter_004:in_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                      : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_002:src1_data -> width_adapter_004:in_data
	signal rsp_xbar_demux_002_src1_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_002:src1_channel -> width_adapter_004:in_channel
	signal rsp_xbar_demux_002_src1_ready                                                                     : std_logic;                      -- width_adapter_004:in_ready -> rsp_xbar_demux_002:src1_ready
	signal width_adapter_004_src_endofpacket                                                                 : std_logic;                      -- width_adapter_004:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal width_adapter_004_src_valid                                                                       : std_logic;                      -- width_adapter_004:out_valid -> rsp_xbar_mux_001:sink2_valid
	signal width_adapter_004_src_startofpacket                                                               : std_logic;                      -- width_adapter_004:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal width_adapter_004_src_data                                                                        : std_logic_vector(114 downto 0); -- width_adapter_004:out_data -> rsp_xbar_mux_001:sink2_data
	signal width_adapter_004_src_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                     : std_logic_vector(3 downto 0);   -- width_adapter_004:out_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src3_endofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src3_endofpacket -> width_adapter_005:in_endofpacket
	signal rsp_xbar_demux_002_src3_valid                                                                     : std_logic;                      -- rsp_xbar_demux_002:src3_valid -> width_adapter_005:in_valid
	signal rsp_xbar_demux_002_src3_startofpacket                                                             : std_logic;                      -- rsp_xbar_demux_002:src3_startofpacket -> width_adapter_005:in_startofpacket
	signal rsp_xbar_demux_002_src3_data                                                                      : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_002:src3_data -> width_adapter_005:in_data
	signal rsp_xbar_demux_002_src3_channel                                                                   : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_002:src3_channel -> width_adapter_005:in_channel
	signal rsp_xbar_demux_002_src3_ready                                                                     : std_logic;                      -- width_adapter_005:in_ready -> rsp_xbar_demux_002:src3_ready
	signal width_adapter_005_src_endofpacket                                                                 : std_logic;                      -- width_adapter_005:out_endofpacket -> vga_m1_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal width_adapter_005_src_valid                                                                       : std_logic;                      -- width_adapter_005:out_valid -> vga_m1_translator_avalon_universal_master_0_agent:rp_valid
	signal width_adapter_005_src_startofpacket                                                               : std_logic;                      -- width_adapter_005:out_startofpacket -> vga_m1_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal width_adapter_005_src_data                                                                        : std_logic_vector(114 downto 0); -- width_adapter_005:out_data -> vga_m1_translator_avalon_universal_master_0_agent:rp_data
	signal width_adapter_005_src_channel                                                                     : std_logic_vector(3 downto 0);   -- width_adapter_005:out_channel -> vga_m1_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_cmd_valid_data                                                                            : std_logic_vector(3 downto 0);   -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                        : std_logic_vector(3 downto 0);   -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal limiter_002_cmd_valid_data                                                                        : std_logic_vector(13 downto 0);  -- limiter_002:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	signal nios2_fast_d_irq_irq                                                                              : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_fast:d_irq
	signal irq_mapper_receiver0_irq                                                                          : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                                                     : std_logic_vector(0 downto 0);   -- systimer:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                                                          : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- sysuart:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver2_irq                                                                          : std_logic;                      -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_002_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver3_irq                                                                          : std_logic;                      -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_003_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- psw:irq -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver4_irq                                                                          : std_logic;                      -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	signal irq_synchronizer_004_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- spu:avs_s1_irq -> irq_synchronizer_004:receiver_irq
	signal irq_mapper_receiver5_irq                                                                          : std_logic;                      -- irq_synchronizer_005:sender_irq -> irq_mapper:receiver5_irq
	signal irq_synchronizer_005_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- ps2_keyboard:irq -> irq_synchronizer_005:receiver_irq
	signal irq_mapper_receiver6_irq                                                                          : std_logic;                      -- irq_synchronizer_006:sender_irq -> irq_mapper:receiver6_irq
	signal irq_synchronizer_006_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- mmcdma:irq -> irq_synchronizer_006:receiver_irq
	signal irq_mapper_receiver7_irq                                                                          : std_logic;                      -- irq_synchronizer_007:sender_irq -> irq_mapper:receiver7_irq
	signal irq_synchronizer_007_receiver_irq                                                                 : std_logic_vector(0 downto 0);   -- vga:irq_s1 -> irq_synchronizer_007:receiver_irq
	signal sys_reset_reset_n_ports_inv                                                                       : std_logic;                      -- sys_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal sdram_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_write:inv -> sdram:az_wr_n
	signal sdram_s1_translator_avalon_anti_slave_0_read_ports_inv                                            : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_read:inv -> sdram:az_rd_n
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                      : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram:az_be_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal sysuart_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                      -- sysuart_s1_translator_avalon_anti_slave_0_write:inv -> sysuart:write_n
	signal sysuart_s1_translator_avalon_anti_slave_0_read_ports_inv                                          : std_logic;                      -- sysuart_s1_translator_avalon_anti_slave_0_read:inv -> sysuart:read_n
	signal systimer_s1_translator_avalon_anti_slave_0_write_ports_inv                                        : std_logic;                      -- systimer_s1_translator_avalon_anti_slave_0_write:inv -> systimer:write_n
	signal led_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                      -- led_s1_translator_avalon_anti_slave_0_write:inv -> led:write_n
	signal led_7seg_s1_translator_avalon_anti_slave_0_write_ports_inv                                        : std_logic;                      -- led_7seg_s1_translator_avalon_anti_slave_0_write:inv -> led_7seg:write_n
	signal psw_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                      -- psw_s1_translator_avalon_anti_slave_0_write:inv -> psw:write_n
	signal gpio1_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                      -- gpio1_s1_translator_avalon_anti_slave_0_write:inv -> gpio1:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                          : std_logic;                      -- rst_controller_reset_out_reset:inv -> [dipsw:reset_n, gpio1:reset_n, jtag_uart:rst_n, led:reset_n, led_7seg:reset_n, psw:reset_n, sysid:reset_n, systimer:reset_n, sysuart:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                                      : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [nios2_fast:reset_n, sdram:reset_n]

begin

	peripherals_bridge : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			ADDRESS_WIDTH       => 14,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk_40mhz_clk,                                                      --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                                     -- m0_reset.reset
			s0_clk           => clk_100mhz_clk,                                                     --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                                 -- s0_reset.reset
			s0_waitrequest   => peripherals_bridge_s0_translator_avalon_anti_slave_0_waitrequest,   --       s0.waitrequest
			s0_readdata      => peripherals_bridge_s0_translator_avalon_anti_slave_0_readdata,      --         .readdata
			s0_readdatavalid => peripherals_bridge_s0_translator_avalon_anti_slave_0_readdatavalid, --         .readdatavalid
			s0_burstcount    => peripherals_bridge_s0_translator_avalon_anti_slave_0_burstcount,    --         .burstcount
			s0_writedata     => peripherals_bridge_s0_translator_avalon_anti_slave_0_writedata,     --         .writedata
			s0_address       => peripherals_bridge_s0_translator_avalon_anti_slave_0_address,       --         .address
			s0_write         => peripherals_bridge_s0_translator_avalon_anti_slave_0_write,         --         .write
			s0_read          => peripherals_bridge_s0_translator_avalon_anti_slave_0_read,          --         .read
			s0_byteenable    => peripherals_bridge_s0_translator_avalon_anti_slave_0_byteenable,    --         .byteenable
			s0_debugaccess   => peripherals_bridge_s0_translator_avalon_anti_slave_0_debugaccess,   --         .debugaccess
			m0_waitrequest   => peripherals_bridge_m0_waitrequest,                                  --       m0.waitrequest
			m0_readdata      => peripherals_bridge_m0_readdata,                                     --         .readdata
			m0_readdatavalid => peripherals_bridge_m0_readdatavalid,                                --         .readdatavalid
			m0_burstcount    => peripherals_bridge_m0_burstcount,                                   --         .burstcount
			m0_writedata     => peripherals_bridge_m0_writedata,                                    --         .writedata
			m0_address       => peripherals_bridge_m0_address,                                      --         .address
			m0_write         => peripherals_bridge_m0_write,                                        --         .write
			m0_read          => peripherals_bridge_m0_read,                                         --         .read
			m0_byteenable    => peripherals_bridge_m0_byteenable,                                   --         .byteenable
			m0_debugaccess   => peripherals_bridge_m0_debugaccess                                   --         .debugaccess
		);

	nios2_fast : component cineraria_core_nios2_fast
		port map (
			clk                                   => clk_100mhz_clk,                                                          --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                            --                   reset_n.reset_n
			d_address                             => nios2_fast_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios2_fast_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios2_fast_data_master_read,                                             --                          .read
			d_readdata                            => nios2_fast_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios2_fast_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios2_fast_data_master_write,                                            --                          .write
			d_writedata                           => nios2_fast_data_master_writedata,                                        --                          .writedata
			d_burstcount                          => nios2_fast_data_master_burstcount,                                       --                          .burstcount
			d_readdatavalid                       => nios2_fast_data_master_readdatavalid,                                    --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios2_fast_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios2_fast_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios2_fast_instruction_master_read,                                      --                          .read
			i_readdata                            => nios2_fast_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios2_fast_instruction_master_waitrequest,                               --                          .waitrequest
			i_burstcount                          => nios2_fast_instruction_master_burstcount,                                --                          .burstcount
			i_readdatavalid                       => nios2_fast_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => nios2_fast_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                                    --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			A_ci_multi_done                       => nios2_fast_custom_instruction_master_done,                               -- custom_instruction_master.done
			A_ci_multi_result                     => nios2_fast_custom_instruction_master_multi_result,                       --                          .multi_result
			A_ci_multi_a                          => nios2_fast_custom_instruction_master_multi_a,                            --                          .multi_a
			A_ci_multi_b                          => nios2_fast_custom_instruction_master_multi_b,                            --                          .multi_b
			A_ci_multi_c                          => nios2_fast_custom_instruction_master_multi_c,                            --                          .multi_c
			A_ci_multi_clk_en                     => nios2_fast_custom_instruction_master_clk_en,                             --                          .clk_en
			A_ci_multi_clock                      => nios2_fast_custom_instruction_master_clk,                                --                          .clk
			A_ci_multi_reset                      => nios2_fast_custom_instruction_master_reset,                              --                          .reset
			A_ci_multi_dataa                      => nios2_fast_custom_instruction_master_multi_dataa,                        --                          .multi_dataa
			A_ci_multi_datab                      => nios2_fast_custom_instruction_master_multi_datab,                        --                          .multi_datab
			A_ci_multi_n                          => nios2_fast_custom_instruction_master_multi_n,                            --                          .multi_n
			A_ci_multi_readra                     => nios2_fast_custom_instruction_master_multi_readra,                       --                          .multi_readra
			A_ci_multi_readrb                     => nios2_fast_custom_instruction_master_multi_readrb,                       --                          .multi_readrb
			A_ci_multi_start                      => nios2_fast_custom_instruction_master_start,                              --                          .start
			A_ci_multi_writerc                    => nios2_fast_custom_instruction_master_multi_writerc                       --                          .multi_writerc
		);

	nios_custom_instr_fpoint : component fpoint_wrapper
		generic map (
			useDivider => 0
		)
		port map (
			clk    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk,    -- s1.clk
			clk_en => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --   .clk_en
			dataa  => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  --   .dataa
			datab  => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --   .datab
			n      => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n,      --   .n
			reset  => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --   .reset
			start  => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start,  --   .start
			done   => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done,   --   .done
			result => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result  --   .result
		);

	jtag_uart : component cineraria_core_jtag_uart
		port map (
			clk            => clk_40mhz_clk,                                                              --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_002_receiver_irq(0)                                        --               irq.irq
		);

	sysuart : component cineraria_core_sysuart
		port map (
			clk           => clk_40mhz_clk,                                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address       => sysuart_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			begintransfer => sysuart_s1_translator_avalon_anti_slave_0_begintransfer,   --                    .begintransfer
			chipselect    => sysuart_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			read_n        => sysuart_s1_translator_avalon_anti_slave_0_read_ports_inv,  --                    .read_n
			write_n       => sysuart_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata     => sysuart_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			readdata      => sysuart_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			dataavailable => open,                                                      --                    .dataavailable
			readyfordata  => open,                                                      --                    .readyfordata
			rxd           => sysuart_rxd,                                               -- external_connection.export
			txd           => sysuart_txd,                                               --                    .export
			cts_n         => sysuart_cts_n,                                             --                    .export
			rts_n         => sysuart_rts_n,                                             --                    .export
			irq           => irq_synchronizer_001_receiver_irq(0)                       --                 irq.irq
		);

	sdram : component cineraria_core_sdram
		port map (
			clk            => clk_100mhz_clk,                                               --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                 -- reset.reset_n
			az_addr        => sdram_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => sdr_addr,                                                     --  wire.export
			zs_ba          => sdr_ba,                                                       --      .export
			zs_cas_n       => sdr_cas_n,                                                    --      .export
			zs_cke         => sdr_cke,                                                      --      .export
			zs_cs_n        => sdr_cs_n,                                                     --      .export
			zs_dq          => sdr_dq,                                                       --      .export
			zs_dqm         => sdr_dqm,                                                      --      .export
			zs_ras_n       => sdr_ras_n,                                                    --      .export
			zs_we_n        => sdr_we_n                                                      --      .export
		);

	ipl_memory : component cineraria_core_ipl_memory
		port map (
			clk        => clk_100mhz_clk,                                          --   clk1.clk
			address    => ipl_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => ipl_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => ipl_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => ipl_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => ipl_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => ipl_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => ipl_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,                      -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req                   --       .reset_req
		);

	sysid : component cineraria_core_sysid
		port map (
			clock    => clk_40mhz_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                      --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	systimer : component cineraria_core_systimer
		port map (
			clk        => clk_40mhz_clk,                                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			address    => systimer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => systimer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => systimer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => systimer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => systimer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_receiver_irq(0)                            --   irq.irq
		);

	led : component cineraria_core_led
		port map (
			clk        => clk_40mhz_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => led_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => led_export                                             -- external_connection.export
		);

	led_7seg : component cineraria_core_led_7seg
		port map (
			clk        => clk_40mhz_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => led_7seg_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_7seg_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_7seg_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_7seg_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_7seg_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => led_7seg_export                                             -- external_connection.export
		);

	psw : component cineraria_core_psw
		port map (
			clk        => clk_40mhz_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => psw_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => psw_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => psw_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => psw_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => psw_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => psw_export,                                            -- external_connection.export
			irq        => irq_synchronizer_003_receiver_irq(0)                   --                 irq.irq
		);

	dipsw : component cineraria_core_dipsw
		port map (
			clk      => clk_40mhz_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address  => dipsw_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => dipsw_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => dipsw_export                                      -- external_connection.export
		);

	nios_custom_instr_pixelsimd : component pixelsimd
		port map (
			dataa  => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa,  -- nios_custom_instruction_slave_0.dataa
			datab  => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab,  --                                .datab
			result => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result, --                                .result
			clk    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk,    --                                .clk
			clk_en => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en, --                                .clk_en
			reset  => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset,  --                                .reset
			start  => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start,  --                                .start
			done   => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done,   --                                .done
			n      => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n       --                                .n
		);

	spu : component avalonif_spu
		port map (
			csi_global_clock     => clk_40mhz_clk,                                     --       global.clk
			csi_global_reset     => rst_controller_reset_out_reset,                    -- global_reset.reset
			csi_m1_clock         => clk_100mhz_clk,                                    --     m1_clock.clk
			avm_m1_address       => spu_m1_address,                                    --           m1.address
			avm_m1_burstcount    => spu_m1_burstcount,                                 --             .burstcount
			avm_m1_read          => spu_m1_read,                                       --             .read
			avm_m1_readdata      => spu_m1_readdata,                                   --             .readdata
			avm_m1_readdatavalid => spu_m1_readdatavalid,                              --             .readdatavalid
			avm_m1_waitrequest   => spu_m1_waitrequest,                                --             .waitrequest
			avs_s1_address       => spu_s1_translator_avalon_anti_slave_0_address,     --           s1.address
			avs_s1_chipselect    => spu_s1_translator_avalon_anti_slave_0_chipselect,  --             .chipselect
			avs_s1_read          => spu_s1_translator_avalon_anti_slave_0_read,        --             .read
			avs_s1_write         => spu_s1_translator_avalon_anti_slave_0_write,       --             .write
			avs_s1_byteenable    => spu_s1_translator_avalon_anti_slave_0_byteenable,  --             .byteenable
			avs_s1_readdata      => spu_s1_translator_avalon_anti_slave_0_readdata,    --             .readdata
			avs_s1_writedata     => spu_s1_translator_avalon_anti_slave_0_writedata,   --             .writedata
			avs_s1_waitrequest   => spu_s1_translator_avalon_anti_slave_0_waitrequest, --             .waitrequest
			avs_s1_irq           => irq_synchronizer_004_receiver_irq(0),              --       irq_s1.irq
			clk_128fs            => spu_clk_128fs,                                     --  conduit_end.export
			DAC_BCLK             => spu_DAC_BCLK,                                      --             .export
			DAC_LRCK             => spu_DAC_LRCK,                                      --             .export
			DAC_DATA             => spu_DAC_DATA,                                      --             .export
			AUD_L                => spu_AUD_L,                                         --             .export
			AUD_R                => spu_AUD_R,                                         --             .export
			SPDIF                => spu_SPDIF                                          --             .export
		);

	mmcdma : component avalonif_mmcdma
		generic map (
			SYSTEMCLOCKINFO => 40000000
		)
		port map (
			clk        => clk_40mhz_clk,                                       --       clock_reset.clk
			reset      => rst_controller_reset_out_reset,                      -- clock_reset_reset.reset
			chipselect => mmcdma_s1_translator_avalon_anti_slave_0_chipselect, --                s1.chipselect
			address    => mmcdma_s1_translator_avalon_anti_slave_0_address,    --                  .address
			read       => mmcdma_s1_translator_avalon_anti_slave_0_read,       --                  .read
			readdata   => mmcdma_s1_translator_avalon_anti_slave_0_readdata,   --                  .readdata
			write      => mmcdma_s1_translator_avalon_anti_slave_0_write,      --                  .write
			writedata  => mmcdma_s1_translator_avalon_anti_slave_0_writedata,  --                  .writedata
			MMC_nCS    => mmc_nCS,                                             --       conduit_end.export
			MMC_SCK    => mmc_SCK,                                             --                  .export
			MMC_SDO    => mmc_SDO,                                             --                  .export
			MMC_SDI    => mmc_SDI,                                             --                  .export
			MMC_CD     => mmc_CD,                                              --                  .export
			MMC_WP     => mmc_WP,                                              --                  .export
			irq        => irq_synchronizer_006_receiver_irq(0)                 --  interrupt_sender.irq
		);

	ps2_keyboard : component ps2_component
		port map (
			clk         => clk_40mhz_clk,                                                        --       clock_reset.clk
			reset       => rst_controller_reset_out_reset,                                       -- clock_reset_reset.reset
			address     => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_address(0),  --      avalon_slave.address
			chipselect  => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_chipselect,  --                  .chipselect
			byteenable  => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_byteenable,  --                  .byteenable
			read        => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_read,        --                  .read
			write       => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_write,       --                  .write
			writedata   => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_writedata,   --                  .writedata
			readdata    => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_readdata,    --                  .readdata
			waitrequest => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_waitrequest, --                  .waitrequest
			PS2_CLK     => ps2kb_CLK,                                                            --       conduit_end.export
			PS2_DAT     => ps2kb_DAT,                                                            --                  .export
			irq         => irq_synchronizer_005_receiver_irq(0)                                  --  interrupt_sender.irq
		);

	gpio1 : component cineraria_core_gpio1
		port map (
			clk        => clk_40mhz_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => gpio1_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => gpio1_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => gpio1_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => gpio1_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => gpio1_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			bidir_port => gpio1_export                                             -- external_connection.export
		);

	vga : component vga_component
		generic map (
			LINEOFFSETBYTES => 2048,
			H_TOTAL         => 525,
			H_SYNC          => 40,
			H_BACKP         => 0,
			H_ACTIVE        => 480,
			V_TOTAL         => 288,
			V_SYNC          => 3,
			V_BACKP         => 0,
			V_ACTIVE        => 272
		)
		port map (
			video_clk            => vga_clk,                                         --     ext.export
			video_rout           => vga_rout,                                        --        .export
			video_gout           => vga_gout,                                        --        .export
			video_bout           => vga_bout,                                        --        .export
			video_hsync_n        => vga_hsync_n,                                     --        .export
			video_vsync_n        => vga_vsync_n,                                     --        .export
			video_enable         => vga_enable,                                      --        .export
			avm_m1_address       => vga_m1_address,                                  --      m1.address
			avm_m1_waitrequest   => vga_m1_waitrequest,                              --        .waitrequest
			avm_m1_burstcount    => vga_m1_burstcount,                               --        .burstcount
			avm_m1_read          => vga_m1_read,                                     --        .read
			avm_m1_readdata      => vga_m1_readdata,                                 --        .readdata
			avm_m1_readdatavalid => vga_m1_readdatavalid,                            --        .readdatavalid
			avs_s1_address       => vga_s1_translator_avalon_anti_slave_0_address,   --      s1.address
			avs_s1_read          => vga_s1_translator_avalon_anti_slave_0_read,      --        .read
			avs_s1_readdata      => vga_s1_translator_avalon_anti_slave_0_readdata,  --        .readdata
			avs_s1_write         => vga_s1_translator_avalon_anti_slave_0_write,     --        .write
			avs_s1_writedata     => vga_s1_translator_avalon_anti_slave_0_writedata, --        .writedata
			irq_s1               => irq_synchronizer_007_receiver_irq(0),            --     irq.irq
			s1_clk               => clk_40mhz_clk,                                   --   s_clk.clk
			m1_clk               => clk_100mhz_clk,                                  --   m_clk.clk
			g_reset              => rst_controller_reset_out_reset                   -- g_reset.reset
		);

	blcon : component backlight_control
		port map (
			reset         => rst_controller_reset_out_reset,                    -- reset.reset
			clk           => clk_40mhz_clk,                                     -- clock.clk
			readdata      => blcon_s1_translator_avalon_anti_slave_0_readdata,  --    s1.readdata
			write         => blcon_s1_translator_avalon_anti_slave_0_write,     --      .write
			writedata     => blcon_s1_translator_avalon_anti_slave_0_writedata, --      .writedata
			read          => blcon_s1_translator_avalon_anti_slave_0_read,      --      .read
			backlight_on  => blcon_on,                                          --   ext.export
			backlight_pwm => blcon_pwm                                          --      .export
		);

	nios2_fast_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 0
		)
		port map (
			ci_slave_result         => open,                                                                    --        ci_slave.result
			ci_slave_multi_clk      => nios2_fast_custom_instruction_master_clk,                                --                .clk
			ci_slave_multi_reset    => nios2_fast_custom_instruction_master_reset,                              --                .reset
			ci_slave_multi_clken    => nios2_fast_custom_instruction_master_clk_en,                             --                .clk_en
			ci_slave_multi_start    => nios2_fast_custom_instruction_master_start,                              --                .start
			ci_slave_multi_done     => nios2_fast_custom_instruction_master_done,                               --                .done
			ci_slave_multi_dataa    => nios2_fast_custom_instruction_master_multi_dataa,                        --                .multi_dataa
			ci_slave_multi_datab    => nios2_fast_custom_instruction_master_multi_datab,                        --                .multi_datab
			ci_slave_multi_result   => nios2_fast_custom_instruction_master_multi_result,                       --                .multi_result
			ci_slave_multi_n        => nios2_fast_custom_instruction_master_multi_n,                            --                .multi_n
			ci_slave_multi_readra   => nios2_fast_custom_instruction_master_multi_readra,                       --                .multi_readra
			ci_slave_multi_readrb   => nios2_fast_custom_instruction_master_multi_readrb,                       --                .multi_readrb
			ci_slave_multi_writerc  => nios2_fast_custom_instruction_master_multi_writerc,                      --                .multi_writerc
			ci_slave_multi_a        => nios2_fast_custom_instruction_master_multi_a,                            --                .multi_a
			ci_slave_multi_b        => nios2_fast_custom_instruction_master_multi_b,                            --                .multi_b
			ci_slave_multi_c        => nios2_fast_custom_instruction_master_multi_c,                            --                .multi_c
			comb_ci_master_result   => open,                                                                    --  comb_ci_master.result
			multi_ci_master_clk     => nios2_fast_custom_instruction_master_translator_multi_ci_master_clk,     -- multi_ci_master.clk
			multi_ci_master_reset   => nios2_fast_custom_instruction_master_translator_multi_ci_master_reset,   --                .reset
			multi_ci_master_clken   => nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en,  --                .clk_en
			multi_ci_master_start   => nios2_fast_custom_instruction_master_translator_multi_ci_master_start,   --                .start
			multi_ci_master_done    => nios2_fast_custom_instruction_master_translator_multi_ci_master_done,    --                .done
			multi_ci_master_dataa   => nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa,   --                .dataa
			multi_ci_master_datab   => nios2_fast_custom_instruction_master_translator_multi_ci_master_datab,   --                .datab
			multi_ci_master_result  => nios2_fast_custom_instruction_master_translator_multi_ci_master_result,  --                .result
			multi_ci_master_n       => nios2_fast_custom_instruction_master_translator_multi_ci_master_n,       --                .n
			multi_ci_master_readra  => nios2_fast_custom_instruction_master_translator_multi_ci_master_readra,  --                .readra
			multi_ci_master_readrb  => nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb,  --                .readrb
			multi_ci_master_writerc => nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc, --                .writerc
			multi_ci_master_a       => nios2_fast_custom_instruction_master_translator_multi_ci_master_a,       --                .a
			multi_ci_master_b       => nios2_fast_custom_instruction_master_translator_multi_ci_master_b,       --                .b
			multi_ci_master_c       => nios2_fast_custom_instruction_master_translator_multi_ci_master_c,       --                .c
			ci_slave_dataa          => "00000000000000000000000000000000",                                      --     (terminated)
			ci_slave_datab          => "00000000000000000000000000000000",                                      --     (terminated)
			ci_slave_n              => "00000000",                                                              --     (terminated)
			ci_slave_readra         => '0',                                                                     --     (terminated)
			ci_slave_readrb         => '0',                                                                     --     (terminated)
			ci_slave_writerc        => '0',                                                                     --     (terminated)
			ci_slave_a              => "00000",                                                                 --     (terminated)
			ci_slave_b              => "00000",                                                                 --     (terminated)
			ci_slave_c              => "00000",                                                                 --     (terminated)
			ci_slave_ipending       => "00000000000000000000000000000000",                                      --     (terminated)
			ci_slave_estatus        => '0',                                                                     --     (terminated)
			comb_ci_master_dataa    => open,                                                                    --     (terminated)
			comb_ci_master_datab    => open,                                                                    --     (terminated)
			comb_ci_master_n        => open,                                                                    --     (terminated)
			comb_ci_master_readra   => open,                                                                    --     (terminated)
			comb_ci_master_readrb   => open,                                                                    --     (terminated)
			comb_ci_master_writerc  => open,                                                                    --     (terminated)
			comb_ci_master_a        => open,                                                                    --     (terminated)
			comb_ci_master_b        => open,                                                                    --     (terminated)
			comb_ci_master_c        => open,                                                                    --     (terminated)
			comb_ci_master_ipending => open,                                                                    --     (terminated)
			comb_ci_master_estatus  => open                                                                     --     (terminated)
		);

	nios2_fast_custom_instruction_master_multi_xconnect : component cineraria_core_nios2_fast_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa      => nios2_fast_custom_instruction_master_translator_multi_ci_master_dataa,   --   ci_slave.dataa
			ci_slave_datab      => nios2_fast_custom_instruction_master_translator_multi_ci_master_datab,   --           .datab
			ci_slave_result     => nios2_fast_custom_instruction_master_translator_multi_ci_master_result,  --           .result
			ci_slave_n          => nios2_fast_custom_instruction_master_translator_multi_ci_master_n,       --           .n
			ci_slave_readra     => nios2_fast_custom_instruction_master_translator_multi_ci_master_readra,  --           .readra
			ci_slave_readrb     => nios2_fast_custom_instruction_master_translator_multi_ci_master_readrb,  --           .readrb
			ci_slave_writerc    => nios2_fast_custom_instruction_master_translator_multi_ci_master_writerc, --           .writerc
			ci_slave_a          => nios2_fast_custom_instruction_master_translator_multi_ci_master_a,       --           .a
			ci_slave_b          => nios2_fast_custom_instruction_master_translator_multi_ci_master_b,       --           .b
			ci_slave_c          => nios2_fast_custom_instruction_master_translator_multi_ci_master_c,       --           .c
			ci_slave_ipending   => open,                                                                    --           .ipending
			ci_slave_estatus    => open,                                                                    --           .estatus
			ci_slave_clk        => nios2_fast_custom_instruction_master_translator_multi_ci_master_clk,     --           .clk
			ci_slave_reset      => nios2_fast_custom_instruction_master_translator_multi_ci_master_reset,   --           .reset
			ci_slave_clken      => nios2_fast_custom_instruction_master_translator_multi_ci_master_clk_en,  --           .clk_en
			ci_slave_start      => nios2_fast_custom_instruction_master_translator_multi_ci_master_start,   --           .start
			ci_slave_done       => nios2_fast_custom_instruction_master_translator_multi_ci_master_done,    --           .done
			ci_master0_dataa    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa,    -- ci_master0.dataa
			ci_master0_datab    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab,    --           .datab
			ci_master0_result   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result,   --           .result
			ci_master0_n        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n,        --           .n
			ci_master0_readra   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra,   --           .readra
			ci_master0_readrb   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb,   --           .readrb
			ci_master0_writerc  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc,  --           .writerc
			ci_master0_a        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a,        --           .a
			ci_master0_b        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b,        --           .b
			ci_master0_c        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c,        --           .c
			ci_master0_ipending => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending, --           .ipending
			ci_master0_estatus  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus,  --           .estatus
			ci_master0_clk      => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk,      --           .clk
			ci_master0_reset    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset,    --           .reset
			ci_master0_clken    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en,   --           .clk_en
			ci_master0_start    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start,    --           .start
			ci_master0_done     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done,     --           .done
			ci_master1_dataa    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa,    -- ci_master1.dataa
			ci_master1_datab    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab,    --           .datab
			ci_master1_result   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result,   --           .result
			ci_master1_n        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n,        --           .n
			ci_master1_readra   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra,   --           .readra
			ci_master1_readrb   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb,   --           .readrb
			ci_master1_writerc  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc,  --           .writerc
			ci_master1_a        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a,        --           .a
			ci_master1_b        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b,        --           .b
			ci_master1_c        => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c,        --           .c
			ci_master1_ipending => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending, --           .ipending
			ci_master1_estatus  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus,  --           .estatus
			ci_master1_clk      => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk,      --           .clk
			ci_master1_reset    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset,    --           .reset
			ci_master1_clken    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en,   --           .clk_en
			ci_master1_start    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start,    --           .start
			ci_master1_done     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done      --           .done
		);

	nios2_fast_custom_instruction_master_multi_slave_translator0 : component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator0
		generic map (
			N_WIDTH          => 2,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk       => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done      => nios2_fast_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result   => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_n        => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_n,      --          .n
			ci_master_clk      => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_clk_en, --          .clk_en
			ci_master_reset    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start    => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done     => nios2_fast_custom_instruction_master_multi_slave_translator0_ci_master_done,   --          .done
			ci_master_readra   => open,                                                                          -- (terminated)
			ci_master_readrb   => open,                                                                          -- (terminated)
			ci_master_writerc  => open,                                                                          -- (terminated)
			ci_master_a        => open,                                                                          -- (terminated)
			ci_master_b        => open,                                                                          -- (terminated)
			ci_master_c        => open,                                                                          -- (terminated)
			ci_master_ipending => open,                                                                          -- (terminated)
			ci_master_estatus  => open                                                                           -- (terminated)
		);

	nios2_fast_custom_instruction_master_multi_slave_translator1 : component cineraria_core_nios2_fast_custom_instruction_master_multi_slave_translator1
		generic map (
			N_WIDTH          => 3,
			USE_DONE         => 1,
			NUM_FIXED_CYCLES => 0
		)
		port map (
			ci_slave_dataa     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_dataa,          --  ci_slave.dataa
			ci_slave_datab     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_datab,          --          .datab
			ci_slave_result    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_result,         --          .result
			ci_slave_n         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_n,              --          .n
			ci_slave_readra    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readra,         --          .readra
			ci_slave_readrb    => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_readrb,         --          .readrb
			ci_slave_writerc   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_writerc,        --          .writerc
			ci_slave_a         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_a,              --          .a
			ci_slave_b         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_b,              --          .b
			ci_slave_c         => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_c,              --          .c
			ci_slave_ipending  => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_ipending,       --          .ipending
			ci_slave_estatus   => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_estatus,        --          .estatus
			ci_slave_clk       => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk,            --          .clk
			ci_slave_clken     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_clk_en,         --          .clk_en
			ci_slave_reset     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_reset,          --          .reset
			ci_slave_start     => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_start,          --          .start
			ci_slave_done      => nios2_fast_custom_instruction_master_multi_xconnect_ci_master1_done,           --          .done
			ci_master_dataa    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_datab,  --          .datab
			ci_master_result   => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_result, --          .result
			ci_master_n        => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_n,      --          .n
			ci_master_clk      => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk,    --          .clk
			ci_master_clken    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_clk_en, --          .clk_en
			ci_master_reset    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_reset,  --          .reset
			ci_master_start    => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_start,  --          .start
			ci_master_done     => nios2_fast_custom_instruction_master_multi_slave_translator1_ci_master_done,   --          .done
			ci_master_readra   => open,                                                                          -- (terminated)
			ci_master_readrb   => open,                                                                          -- (terminated)
			ci_master_writerc  => open,                                                                          -- (terminated)
			ci_master_a        => open,                                                                          -- (terminated)
			ci_master_b        => open,                                                                          -- (terminated)
			ci_master_c        => open,                                                                          -- (terminated)
			ci_master_ipending => open,                                                                          -- (terminated)
			ci_master_estatus  => open                                                                           -- (terminated)
		);

	nios2_fast_instruction_master_translator : component cineraria_core_nios2_fast_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 28,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 4,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 6,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 1,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                               --                     reset.reset
			uav_address              => nios2_fast_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_fast_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_fast_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_fast_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_fast_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_fast_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_fast_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_fast_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_fast_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_fast_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_fast_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_fast_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_fast_instruction_master_waitrequest,                                        --                          .waitrequest
			av_burstcount            => nios2_fast_instruction_master_burstcount,                                         --                          .burstcount
			av_read                  => nios2_fast_instruction_master_read,                                               --                          .read
			av_readdata              => nios2_fast_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => nios2_fast_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_byteenable            => "1111",                                                                           --               (terminated)
			av_beginbursttransfer    => '0',                                                                              --               (terminated)
			av_begintransfer         => '0',                                                                              --               (terminated)
			av_chipselect            => '0',                                                                              --               (terminated)
			av_write                 => '0',                                                                              --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                               --               (terminated)
			av_lock                  => '0',                                                                              --               (terminated)
			av_debugaccess           => '0',                                                                              --               (terminated)
			uav_clken                => open,                                                                             --               (terminated)
			av_clken                 => '1',                                                                              --               (terminated)
			uav_response             => "00",                                                                             --               (terminated)
			av_response              => open,                                                                             --               (terminated)
			uav_writeresponserequest => open,                                                                             --               (terminated)
			uav_writeresponsevalid   => '0',                                                                              --               (terminated)
			av_writeresponserequest  => '0',                                                                              --               (terminated)
			av_writeresponsevalid    => open                                                                              --               (terminated)
		);

	nios2_fast_data_master_translator : component cineraria_core_nios2_fast_data_master_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 4,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 6,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 1,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                            --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                        --                     reset.reset
			uav_address              => nios2_fast_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_fast_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_fast_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_fast_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_fast_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_fast_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_fast_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_fast_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_fast_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_fast_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_fast_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_fast_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_fast_data_master_waitrequest,                                        --                          .waitrequest
			av_burstcount            => nios2_fast_data_master_burstcount,                                         --                          .burstcount
			av_byteenable            => nios2_fast_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios2_fast_data_master_read,                                               --                          .read
			av_readdata              => nios2_fast_data_master_readdata,                                           --                          .readdata
			av_readdatavalid         => nios2_fast_data_master_readdatavalid,                                      --                          .readdatavalid
			av_write                 => nios2_fast_data_master_write,                                              --                          .write
			av_writedata             => nios2_fast_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios2_fast_data_master_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	spu_m1_translator : component cineraria_core_spu_m1_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 16,
			AV_BURSTCOUNT_W             => 3,
			AV_BYTEENABLE_W             => 2,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 4,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 2,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 1,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                            --                       clk.clk
			reset                    => rst_controller_002_reset_out_reset,                        --                     reset.reset
			uav_address              => spu_m1_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => spu_m1_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => spu_m1_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => spu_m1_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => spu_m1_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => spu_m1_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => spu_m1_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => spu_m1_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => spu_m1_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => spu_m1_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => spu_m1_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => spu_m1_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => spu_m1_waitrequest,                                        --                          .waitrequest
			av_burstcount            => spu_m1_burstcount,                                         --                          .burstcount
			av_read                  => spu_m1_read,                                               --                          .read
			av_readdata              => spu_m1_readdata,                                           --                          .readdata
			av_readdatavalid         => spu_m1_readdatavalid,                                      --                          .readdatavalid
			av_byteenable            => "11",                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                       --               (terminated)
			av_begintransfer         => '0',                                                       --               (terminated)
			av_chipselect            => '0',                                                       --               (terminated)
			av_write                 => '0',                                                       --               (terminated)
			av_writedata             => "0000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                       --               (terminated)
			av_debugaccess           => '0',                                                       --               (terminated)
			uav_clken                => open,                                                      --               (terminated)
			av_clken                 => '1',                                                       --               (terminated)
			uav_response             => "00",                                                      --               (terminated)
			av_response              => open,                                                      --               (terminated)
			uav_writeresponserequest => open,                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                       --               (terminated)
			av_writeresponsevalid    => open                                                       --               (terminated)
		);

	vga_m1_translator : component cineraria_core_vga_m1_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 10,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 12,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 1,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                            --                       clk.clk
			reset                    => rst_controller_002_reset_out_reset,                        --                     reset.reset
			uav_address              => vga_m1_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => vga_m1_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => vga_m1_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => vga_m1_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => vga_m1_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => vga_m1_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => vga_m1_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => vga_m1_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => vga_m1_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => vga_m1_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => vga_m1_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => vga_m1_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => vga_m1_waitrequest,                                        --                          .waitrequest
			av_burstcount            => vga_m1_burstcount,                                         --                          .burstcount
			av_read                  => vga_m1_read,                                               --                          .read
			av_readdata              => vga_m1_readdata,                                           --                          .readdata
			av_readdatavalid         => vga_m1_readdatavalid,                                      --                          .readdatavalid
			av_byteenable            => "1111",                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                       --               (terminated)
			av_begintransfer         => '0',                                                       --               (terminated)
			av_chipselect            => '0',                                                       --               (terminated)
			av_write                 => '0',                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                        --               (terminated)
			av_lock                  => '0',                                                       --               (terminated)
			av_debugaccess           => '0',                                                       --               (terminated)
			uav_clken                => open,                                                      --               (terminated)
			av_clken                 => '1',                                                       --               (terminated)
			uav_response             => "00",                                                      --               (terminated)
			av_response              => open,                                                      --               (terminated)
			uav_writeresponserequest => open,                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                       --               (terminated)
			av_writeresponsevalid    => open                                                       --               (terminated)
		);

	nios2_fast_jtag_debug_module_translator : component cineraria_core_nios2_fast_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                      --                    reset.reset
			uav_address              => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios2_fast_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                                    --              (terminated)
			av_burstcount            => open,                                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                                    --              (terminated)
			av_lock                  => open,                                                                                    --              (terminated)
			av_chipselect            => open,                                                                                    --              (terminated)
			av_clken                 => open,                                                                                    --              (terminated)
			uav_clken                => '0',                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                    --              (terminated)
			uav_response             => open,                                                                                    --              (terminated)
			av_response              => "00",                                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                                      --              (terminated)
		);

	ipl_memory_s1_translator : component cineraria_core_ipl_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 11,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                    reset.reset
			uav_address              => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ipl_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ipl_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => ipl_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ipl_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => ipl_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => ipl_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => ipl_memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	sdram_s1_translator : component cineraria_core_sdram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                      --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                  --                    reset.reset
			uav_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	peripherals_bridge_s0_translator : component cineraria_core_peripherals_bridge_s0_translator
		generic map (
			AV_ADDRESS_W                   => 14,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100mhz_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                               --                    reset.reset
			uav_address              => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => peripherals_bridge_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => peripherals_bridge_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => peripherals_bridge_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => peripherals_bridge_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => peripherals_bridge_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => peripherals_bridge_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => peripherals_bridge_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => peripherals_bridge_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => peripherals_bridge_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => peripherals_bridge_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	peripherals_bridge_m0_translator : component cineraria_core_peripherals_bridge_m0_translator
		generic map (
			AV_ADDRESS_W                => 14,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 14,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                     reset.reset
			uav_address              => peripherals_bridge_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => peripherals_bridge_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => peripherals_bridge_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => peripherals_bridge_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => peripherals_bridge_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => peripherals_bridge_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => peripherals_bridge_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => peripherals_bridge_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => peripherals_bridge_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => peripherals_bridge_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => peripherals_bridge_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => peripherals_bridge_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => peripherals_bridge_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => peripherals_bridge_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => peripherals_bridge_m0_byteenable,                                         --                          .byteenable
			av_read                  => peripherals_bridge_m0_read,                                               --                          .read
			av_readdata              => peripherals_bridge_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => peripherals_bridge_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => peripherals_bridge_m0_write,                                              --                          .write
			av_writedata             => peripherals_bridge_m0_writedata,                                          --                          .writedata
			av_debugaccess           => peripherals_bridge_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                      --               (terminated)
			av_begintransfer         => '0',                                                                      --               (terminated)
			av_chipselect            => '0',                                                                      --               (terminated)
			av_lock                  => '0',                                                                      --               (terminated)
			uav_clken                => open,                                                                     --               (terminated)
			av_clken                 => '1',                                                                      --               (terminated)
			uav_response             => "00",                                                                     --               (terminated)
			av_response              => open,                                                                     --               (terminated)
			uav_writeresponserequest => open,                                                                     --               (terminated)
			uav_writeresponsevalid   => '0',                                                                      --               (terminated)
			av_writeresponserequest  => '0',                                                                      --               (terminated)
			av_writeresponsevalid    => open                                                                      --               (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component cineraria_core_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	sysuart_s1_translator : component cineraria_core_sysuart_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysuart_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sysuart_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sysuart_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sysuart_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sysuart_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => sysuart_s1_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_chipselect            => sysuart_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	sysid_control_slave_translator : component cineraria_core_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	systimer_s1_translator : component cineraria_core_systimer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => systimer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => systimer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => systimer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => systimer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => systimer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => systimer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => systimer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => systimer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	led_s1_translator : component cineraria_core_led_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => led_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	led_7seg_s1_translator : component cineraria_core_led_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_7seg_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_7seg_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_7seg_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_7seg_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_7seg_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	psw_s1_translator : component cineraria_core_led_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => psw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => psw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => psw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => psw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => psw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => psw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => psw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => psw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => psw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => psw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => psw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => psw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => psw_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => psw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => psw_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => psw_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	dipsw_s1_translator : component cineraria_core_dipsw_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dipsw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => dipsw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                --              (terminated)
			av_read                  => open,                                                                --              (terminated)
			av_writedata             => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_chipselect            => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	spu_s1_translator : component cineraria_core_spu_s1_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => spu_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => spu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => spu_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => spu_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => spu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => spu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => spu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => spu_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => spu_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => spu_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => spu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => spu_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => spu_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => spu_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => spu_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => spu_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => spu_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => spu_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => spu_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	mmcdma_s1_translator : component cineraria_core_mmcdma_s1_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 2,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => mmcdma_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => mmcdma_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => mmcdma_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => mmcdma_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => mmcdma_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => mmcdma_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	ps2_keyboard_avalon_slave_translator : component cineraria_core_ps2_keyboard_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                       --                    reset.reset
			uav_address              => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => ps2_keyboard_avalon_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                                 --              (terminated)
			av_burstcount            => open,                                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                                 --              (terminated)
			av_lock                  => open,                                                                                 --              (terminated)
			av_clken                 => open,                                                                                 --              (terminated)
			uav_clken                => '0',                                                                                  --              (terminated)
			av_debugaccess           => open,                                                                                 --              (terminated)
			av_outputenable          => open,                                                                                 --              (terminated)
			uav_response             => open,                                                                                 --              (terminated)
			av_response              => "00",                                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                                   --              (terminated)
		);

	gpio1_s1_translator : component cineraria_core_led_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => gpio1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => gpio1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => gpio1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => gpio1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => gpio1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	vga_s1_translator : component cineraria_core_vga_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => vga_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => vga_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => vga_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => vga_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => vga_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => vga_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => vga_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => vga_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => vga_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => vga_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => vga_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => vga_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => vga_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => vga_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => vga_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => vga_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_chipselect            => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	blcon_s1_translator : component cineraria_core_blcon_s1_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_40mhz_clk,                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => blcon_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => blcon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => blcon_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => blcon_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => blcon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => blcon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => blcon_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => blcon_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => blcon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_write                 => blcon_s1_translator_avalon_anti_slave_0_write,                       --      avalon_anti_slave_0.write
			av_read                  => blcon_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => blcon_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => blcon_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_address               => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_chipselect            => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	nios2_fast_instruction_master_translator_avalon_universal_master_0_agent : component cineraria_core_nios2_fast_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_BEGIN_BURST           => 99,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_THREAD_ID_H           => 105,
			PKT_THREAD_ID_L           => 105,
			PKT_CACHE_H               => 112,
			PKT_CACHE_L               => 109,
			PKT_DATA_SIDEBAND_H       => 98,
			PKT_DATA_SIDEBAND_L       => 98,
			PKT_QOS_H                 => 100,
			PKT_QOS_L                 => 100,
			PKT_ADDR_SIDEBAND_H       => 97,
			PKT_ADDR_SIDEBAND_L       => 97,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 6,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 31,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                            --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                        -- clk_reset.reset
			av_address              => nios2_fast_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_fast_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_fast_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_fast_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_fast_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_fast_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_fast_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_fast_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_fast_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_fast_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_fast_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                                     --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                                      --          .data
			rp_channel              => limiter_rsp_src_channel,                                                                   --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                             --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                               --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                                     --          .ready
			av_response             => open,                                                                                      -- (terminated)
			av_writeresponserequest => '0',                                                                                       -- (terminated)
			av_writeresponsevalid   => open                                                                                       -- (terminated)
		);

	nios2_fast_data_master_translator_avalon_universal_master_0_agent : component cineraria_core_nios2_fast_instruction_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_BEGIN_BURST           => 99,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_THREAD_ID_H           => 105,
			PKT_THREAD_ID_L           => 105,
			PKT_CACHE_H               => 112,
			PKT_CACHE_L               => 109,
			PKT_DATA_SIDEBAND_H       => 98,
			PKT_DATA_SIDEBAND_L       => 98,
			PKT_QOS_H                 => 100,
			PKT_QOS_L                 => 100,
			PKT_ADDR_SIDEBAND_H       => 97,
			PKT_ADDR_SIDEBAND_L       => 97,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 6,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 63,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                     --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			av_address              => nios2_fast_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_fast_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_fast_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_fast_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_fast_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_fast_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_fast_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_fast_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_fast_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_fast_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_fast_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_001_rsp_src_valid,                                                          --        rp.valid
			rp_data                 => limiter_001_rsp_src_data,                                                           --          .data
			rp_channel              => limiter_001_rsp_src_channel,                                                        --          .channel
			rp_startofpacket        => limiter_001_rsp_src_startofpacket,                                                  --          .startofpacket
			rp_endofpacket          => limiter_001_rsp_src_endofpacket,                                                    --          .endofpacket
			rp_ready                => limiter_001_rsp_src_ready,                                                          --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	spu_m1_translator_avalon_universal_master_0_agent : component cineraria_core_spu_m1_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 90,
			PKT_PROTECTION_L          => 88,
			PKT_BEGIN_BURST           => 81,
			PKT_BURSTWRAP_H           => 73,
			PKT_BURSTWRAP_L           => 68,
			PKT_BURST_SIZE_H          => 76,
			PKT_BURST_SIZE_L          => 74,
			PKT_BURST_TYPE_H          => 78,
			PKT_BURST_TYPE_L          => 77,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_SRC_ID_H              => 84,
			PKT_SRC_ID_L              => 83,
			PKT_DEST_ID_H             => 86,
			PKT_DEST_ID_L             => 85,
			PKT_THREAD_ID_H           => 87,
			PKT_THREAD_ID_L           => 87,
			PKT_CACHE_H               => 94,
			PKT_CACHE_L               => 91,
			PKT_DATA_SIDEBAND_H       => 80,
			PKT_DATA_SIDEBAND_L       => 80,
			PKT_QOS_H                 => 82,
			PKT_QOS_L                 => 82,
			PKT_ADDR_SIDEBAND_H       => 79,
			PKT_ADDR_SIDEBAND_L       => 79,
			PKT_RESPONSE_STATUS_H     => 96,
			PKT_RESPONSE_STATUS_L     => 95,
			ST_DATA_W                 => 97,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 4,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 2,
			BURSTWRAP_VALUE           => 63,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                     --       clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                 -- clk_reset.reset
			av_address              => spu_m1_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => spu_m1_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => spu_m1_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => spu_m1_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => spu_m1_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => spu_m1_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => spu_m1_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => spu_m1_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => spu_m1_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => spu_m1_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => spu_m1_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => spu_m1_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => spu_m1_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => spu_m1_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => spu_m1_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => spu_m1_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_002_src2_valid,                                      --        rp.valid
			rp_data                 => rsp_xbar_demux_002_src2_data,                                       --          .data
			rp_channel              => rsp_xbar_demux_002_src2_channel,                                    --          .channel
			rp_startofpacket        => rsp_xbar_demux_002_src2_startofpacket,                              --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_002_src2_endofpacket,                                --          .endofpacket
			rp_ready                => rsp_xbar_demux_002_src2_ready,                                      --          .ready
			av_response             => open,                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                -- (terminated)
		);

	vga_m1_translator_avalon_universal_master_0_agent : component cineraria_core_vga_m1_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_BEGIN_BURST           => 99,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_THREAD_ID_H           => 105,
			PKT_THREAD_ID_L           => 105,
			PKT_CACHE_H               => 112,
			PKT_CACHE_L               => 109,
			PKT_DATA_SIDEBAND_H       => 98,
			PKT_DATA_SIDEBAND_L       => 98,
			PKT_QOS_H                 => 100,
			PKT_QOS_L                 => 100,
			PKT_ADDR_SIDEBAND_H       => 97,
			PKT_ADDR_SIDEBAND_L       => 97,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 12,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 3,
			BURSTWRAP_VALUE           => 63,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                     --       clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                 -- clk_reset.reset
			av_address              => vga_m1_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => vga_m1_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => vga_m1_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => vga_m1_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => vga_m1_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => vga_m1_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => vga_m1_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => vga_m1_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => vga_m1_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => vga_m1_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => vga_m1_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => vga_m1_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => vga_m1_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => vga_m1_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => vga_m1_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => vga_m1_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => width_adapter_005_src_valid,                                        --        rp.valid
			rp_data                 => width_adapter_005_src_data,                                         --          .data
			rp_channel              => width_adapter_005_src_channel,                                      --          .channel
			rp_startofpacket        => width_adapter_005_src_startofpacket,                                --          .startofpacket
			rp_endofpacket          => width_adapter_005_src_endofpacket,                                  --          .endofpacket
			rp_ready                => width_adapter_005_src_ready,                                        --          .ready
			av_response             => open,                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                -- (terminated)
		);

	nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 99,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 115,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                --       clk_reset.reset
			m0_address              => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                       --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                       --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                        --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                                 --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                     --                .channel
			rf_sink_ready           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                --     (terminated)
		);

	nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 116,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                -- clk_reset.reset
			in_data           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                              -- (terminated)
			csr_read          => '0',                                                                                               -- (terminated)
			csr_write         => '0',                                                                                               -- (terminated)
			csr_readdata      => open,                                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                -- (terminated)
			almost_full_data  => open,                                                                                              -- (terminated)
			almost_empty_data => open,                                                                                              -- (terminated)
			in_empty          => '0',                                                                                               -- (terminated)
			out_empty         => open,                                                                                              -- (terminated)
			in_error          => '0',                                                                                               -- (terminated)
			out_error         => open,                                                                                              -- (terminated)
			in_channel        => '0',                                                                                               -- (terminated)
			out_channel       => open                                                                                               -- (terminated)
		);

	nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                              --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_startofpacket  => '0',                                                                                         -- (terminated)
			in_endofpacket    => '0',                                                                                         -- (terminated)
			out_startofpacket => open,                                                                                        -- (terminated)
			out_endofpacket   => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	ipl_memory_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 99,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 115,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ipl_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                    --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                    --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                     --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                              --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                  --                .channel
			rf_sink_ready           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 116,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                               --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_startofpacket  => '0',                                                                          -- (terminated)
			in_endofpacket    => '0',                                                                          -- (terminated)
			out_startofpacket => open,                                                                         -- (terminated)
			out_endofpacket   => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 81,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 84,
			PKT_SRC_ID_L              => 83,
			PKT_DEST_ID_H             => 86,
			PKT_DEST_ID_L             => 85,
			PKT_BURSTWRAP_H           => 73,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 90,
			PKT_PROTECTION_L          => 88,
			PKT_RESPONSE_STATUS_H     => 96,
			PKT_RESPONSE_STATUS_L     => 95,
			PKT_BURST_SIZE_H          => 76,
			PKT_BURST_SIZE_L          => 74,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 97,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                            --       clk_reset.reset
			m0_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_002_source0_ready,                                               --              cp.ready
			cp_valid                => burst_adapter_002_source0_valid,                                               --                .valid
			cp_data                 => burst_adapter_002_source0_data,                                                --                .data
			cp_startofpacket        => burst_adapter_002_source0_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => burst_adapter_002_source0_endofpacket,                                         --                .endofpacket
			cp_channel              => burst_adapter_002_source0_channel,                                             --                .channel
			rf_sink_ready           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 98,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component cineraria_core_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                      -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                    -- (terminated)
			csr_read          => '0',                                                                     -- (terminated)
			csr_write         => '0',                                                                     -- (terminated)
			csr_readdata      => open,                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                      -- (terminated)
			almost_full_data  => open,                                                                    -- (terminated)
			almost_empty_data => open,                                                                    -- (terminated)
			in_startofpacket  => '0',                                                                     -- (terminated)
			in_endofpacket    => '0',                                                                     -- (terminated)
			out_startofpacket => open,                                                                    -- (terminated)
			out_endofpacket   => open,                                                                    -- (terminated)
			in_empty          => '0',                                                                     -- (terminated)
			out_empty         => open,                                                                    -- (terminated)
			in_error          => '0',                                                                     -- (terminated)
			out_error         => open,                                                                    -- (terminated)
			in_channel        => '0',                                                                     -- (terminated)
			out_channel       => open                                                                     -- (terminated)
		);

	peripherals_bridge_s0_translator_avalon_universal_slave_0_agent : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 99,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 102,
			PKT_SRC_ID_L              => 101,
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 108,
			PKT_PROTECTION_L          => 106,
			PKT_RESPONSE_STATUS_H     => 114,
			PKT_RESPONSE_STATUS_L     => 113,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 115,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100mhz_clk,                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_003_source0_ready,                                                            --              cp.ready
			cp_valid                => burst_adapter_003_source0_valid,                                                            --                .valid
			cp_data                 => burst_adapter_003_source0_data,                                                             --                .data
			cp_startofpacket        => burst_adapter_003_source0_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => burst_adapter_003_source0_endofpacket,                                                      --                .endofpacket
			cp_channel              => burst_adapter_003_source0_channel,                                                          --                .channel
			rf_sink_ready           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 116,
			FIFO_DEPTH          => 9,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo : component cineraria_core_nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 16,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100mhz_clk,                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                 -- (terminated)
			csr_read          => '0',                                                                                  -- (terminated)
			csr_write         => '0',                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                   -- (terminated)
			almost_full_data  => open,                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                 -- (terminated)
			in_startofpacket  => '0',                                                                                  -- (terminated)
			in_endofpacket    => '0',                                                                                  -- (terminated)
			out_startofpacket => open,                                                                                 -- (terminated)
			out_endofpacket   => open,                                                                                 -- (terminated)
			in_empty          => '0',                                                                                  -- (terminated)
			out_empty         => open,                                                                                 -- (terminated)
			in_error          => '0',                                                                                  -- (terminated)
			out_error         => open,                                                                                 -- (terminated)
			in_channel        => '0',                                                                                  -- (terminated)
			out_channel       => open                                                                                  -- (terminated)
		);

	peripherals_bridge_m0_translator_avalon_universal_master_0_agent : component cineraria_core_peripherals_bridge_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_BEGIN_BURST           => 67,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			PKT_BURST_TYPE_H          => 64,
			PKT_BURST_TYPE_L          => 63,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_THREAD_ID_H           => 77,
			PKT_THREAD_ID_L           => 77,
			PKT_CACHE_H               => 84,
			PKT_CACHE_L               => 81,
			PKT_DATA_SIDEBAND_H       => 66,
			PKT_DATA_SIDEBAND_L       => 66,
			PKT_QOS_H                 => 68,
			PKT_QOS_L                 => 68,
			PKT_ADDR_SIDEBAND_H       => 65,
			PKT_ADDR_SIDEBAND_L       => 65,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			ST_DATA_W                 => 87,
			ST_CHANNEL_W              => 14,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			av_address              => peripherals_bridge_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => peripherals_bridge_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => peripherals_bridge_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => peripherals_bridge_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => peripherals_bridge_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => peripherals_bridge_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => peripherals_bridge_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => peripherals_bridge_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => peripherals_bridge_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => peripherals_bridge_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => peripherals_bridge_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_002_rsp_src_valid,                                                         --        rp.valid
			rp_data                 => limiter_002_rsp_src_data,                                                          --          .data
			rp_channel              => limiter_002_rsp_src_channel,                                                       --          .channel
			rp_startofpacket        => limiter_002_rsp_src_startofpacket,                                                 --          .startofpacket
			rp_endofpacket          => limiter_002_rsp_src_endofpacket,                                                   --          .endofpacket
			rp_ready                => limiter_002_rsp_src_ready,                                                         --          .ready
			av_response             => open,                                                                              -- (terminated)
			av_writeresponserequest => '0',                                                                               -- (terminated)
			av_writeresponsevalid   => open                                                                               -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src0_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src0_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_004_src0_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src0_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src0_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src0_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	sysuart_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysuart_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src1_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src1_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_004_src1_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src1_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src1_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src1_channel,                                                 --                .channel
			rf_sink_ready           => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysuart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysuart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysuart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src2_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src2_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_004_src2_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src2_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src2_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src2_channel,                                                          --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	systimer_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => systimer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => systimer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => systimer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => systimer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src3_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src3_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_004_src3_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src3_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src3_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src3_channel,                                                  --                .channel
			rf_sink_ready           => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	led_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => led_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src4_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src4_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_004_src4_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src4_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src4_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src4_channel,                                             --                .channel
			rf_sink_ready           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			in_data           => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	led_7seg_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_7seg_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src5_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src5_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_004_src5_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src5_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src5_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src5_channel,                                                  --                .channel
			rf_sink_ready           => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_7seg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_7seg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	psw_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => psw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => psw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => psw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => psw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => psw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => psw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => psw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => psw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => psw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => psw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => psw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => psw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => psw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => psw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => psw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => psw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src6_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src6_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_004_src6_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src6_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src6_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src6_channel,                                             --                .channel
			rf_sink_ready           => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => psw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			in_data           => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => psw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => psw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	dipsw_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                 --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dipsw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src7_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src7_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_004_src7_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src7_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src7_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src7_channel,                                               --                .channel
			rf_sink_ready           => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dipsw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dipsw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dipsw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	spu_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => spu_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => spu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => spu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => spu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => spu_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => spu_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => spu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => spu_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => spu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => spu_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => spu_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => spu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => spu_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => spu_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => spu_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => spu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src8_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src8_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_004_src8_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src8_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src8_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src8_channel,                                             --                .channel
			rf_sink_ready           => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => spu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			in_data           => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => spu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => spu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	mmcdma_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => mmcdma_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src9_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src9_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_004_src9_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src9_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src9_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src9_channel,                                                --                .channel
			rf_sink_ready           => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => mmcdma_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => mmcdma_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                 --       clk_reset.reset
			m0_address              => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src10_ready,                                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src10_valid,                                                                 --                .valid
			cp_data                 => cmd_xbar_demux_004_src10_data,                                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src10_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src10_endofpacket,                                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src10_channel,                                                               --                .channel
			rf_sink_ready           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                             --     (terminated)
		);

	ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                 -- clk_reset.reset
			in_data           => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                           -- (terminated)
			csr_read          => '0',                                                                                            -- (terminated)
			csr_write         => '0',                                                                                            -- (terminated)
			csr_readdata      => open,                                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                             -- (terminated)
			almost_full_data  => open,                                                                                           -- (terminated)
			almost_empty_data => open,                                                                                           -- (terminated)
			in_empty          => '0',                                                                                            -- (terminated)
			out_empty         => open,                                                                                           -- (terminated)
			in_error          => '0',                                                                                            -- (terminated)
			out_error         => open,                                                                                           -- (terminated)
			in_channel        => '0',                                                                                            -- (terminated)
			out_channel       => open                                                                                            -- (terminated)
		);

	gpio1_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                 --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => gpio1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src11_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src11_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_004_src11_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src11_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src11_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src11_channel,                                              --                .channel
			rf_sink_ready           => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => gpio1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => gpio1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => gpio1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	vga_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => vga_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => vga_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => vga_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => vga_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => vga_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => vga_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => vga_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => vga_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => vga_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => vga_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => vga_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => vga_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => vga_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => vga_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => vga_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => vga_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src12_ready,                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src12_valid,                                              --                .valid
			cp_data                 => cmd_xbar_demux_004_src12_data,                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src12_startofpacket,                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src12_endofpacket,                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src12_channel,                                            --                .channel
			rf_sink_ready           => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => vga_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			in_data           => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => vga_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => vga_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	blcon_s1_translator_avalon_universal_slave_0_agent : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 67,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 69,
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 59,
			PKT_BURSTWRAP_L           => 59,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 80,
			PKT_PROTECTION_L          => 78,
			PKT_RESPONSE_STATUS_H     => 86,
			PKT_RESPONSE_STATUS_L     => 85,
			PKT_BURST_SIZE_H          => 62,
			PKT_BURST_SIZE_L          => 60,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 87,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_40mhz_clk,                                                                 --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => blcon_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => blcon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => blcon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => blcon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => blcon_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => blcon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => blcon_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => blcon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => blcon_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => blcon_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => blcon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => blcon_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => blcon_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => blcon_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => blcon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_004_src13_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_004_src13_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_004_src13_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_004_src13_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_004_src13_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_004_src13_channel,                                              --                .channel
			rf_sink_ready           => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => blcon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component cineraria_core_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 88,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_40mhz_clk,                                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => blcon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => blcon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	addr_router : component cineraria_core_addr_router
		port map (
			sink_ready         => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_fast_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                     --       src.ready
			src_valid          => addr_router_src_valid,                                                                     --          .valid
			src_data           => addr_router_src_data,                                                                      --          .data
			src_channel        => addr_router_src_channel,                                                                   --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                --          .endofpacket
		);

	addr_router_001 : component cineraria_core_addr_router_001
		port map (
			sink_ready         => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_fast_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                          --       src.ready
			src_valid          => addr_router_001_src_valid,                                                          --          .valid
			src_data           => addr_router_001_src_data,                                                           --          .data
			src_channel        => addr_router_001_src_channel,                                                        --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                     --          .endofpacket
		);

	addr_router_002 : component cineraria_core_addr_router_002
		port map (
			sink_ready         => spu_m1_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => spu_m1_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => spu_m1_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => spu_m1_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => spu_m1_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                 -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                          --       src.ready
			src_valid          => addr_router_002_src_valid,                                          --          .valid
			src_data           => addr_router_002_src_data,                                           --          .data
			src_channel        => addr_router_002_src_channel,                                        --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                  --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                     --          .endofpacket
		);

	addr_router_003 : component cineraria_core_addr_router_003
		port map (
			sink_ready         => vga_m1_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => vga_m1_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => vga_m1_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => vga_m1_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_m1_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                 -- clk_reset.reset
			src_ready          => addr_router_003_src_ready,                                          --       src.ready
			src_valid          => addr_router_003_src_valid,                                          --          .valid
			src_data           => addr_router_003_src_data,                                           --          .data
			src_channel        => addr_router_003_src_channel,                                        --          .channel
			src_startofpacket  => addr_router_003_src_startofpacket,                                  --          .startofpacket
			src_endofpacket    => addr_router_003_src_endofpacket                                     --          .endofpacket
		);

	id_router : component cineraria_core_id_router
		port map (
			sink_ready         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_fast_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                                          --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                     --       src.ready
			src_valid          => id_router_src_valid,                                                                     --          .valid
			src_data           => id_router_src_data,                                                                      --          .data
			src_channel        => id_router_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                --          .endofpacket
		);

	id_router_001 : component cineraria_core_id_router
		port map (
			sink_ready         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ipl_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                  --       src.ready
			src_valid          => id_router_001_src_valid,                                                  --          .valid
			src_data           => id_router_001_src_data,                                                   --          .data
			src_channel        => id_router_001_src_channel,                                                --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                             --          .endofpacket
		);

	id_router_002 : component cineraria_core_id_router_002
		port map (
			sink_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                      --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                  -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                             --       src.ready
			src_valid          => id_router_002_src_valid,                                             --          .valid
			src_data           => id_router_002_src_data,                                              --          .data
			src_channel        => id_router_002_src_channel,                                           --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                        --          .endofpacket
		);

	id_router_003 : component cineraria_core_id_router_003
		port map (
			sink_ready         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => peripherals_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100mhz_clk,                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                          --       src.ready
			src_valid          => id_router_003_src_valid,                                                          --          .valid
			src_data           => id_router_003_src_data,                                                           --          .data
			src_channel        => id_router_003_src_channel,                                                        --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                     --          .endofpacket
		);

	addr_router_004 : component cineraria_core_addr_router_004
		port map (
			sink_ready         => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => peripherals_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => addr_router_004_src_ready,                                                         --       src.ready
			src_valid          => addr_router_004_src_valid,                                                         --          .valid
			src_data           => addr_router_004_src_data,                                                          --          .data
			src_channel        => addr_router_004_src_channel,                                                       --          .channel
			src_startofpacket  => addr_router_004_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => addr_router_004_src_endofpacket                                                    --          .endofpacket
		);

	id_router_004 : component cineraria_core_id_router_004
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                --       src.ready
			src_valid          => id_router_004_src_valid,                                                                --          .valid
			src_data           => id_router_004_src_data,                                                                 --          .data
			src_channel        => id_router_004_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                           --          .endofpacket
		);

	id_router_005 : component cineraria_core_id_router_004
		port map (
			sink_ready         => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysuart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                               --       src.ready
			src_valid          => id_router_005_src_valid,                                               --          .valid
			src_data           => id_router_005_src_data,                                                --          .data
			src_channel        => id_router_005_src_channel,                                             --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                          --          .endofpacket
		);

	id_router_006 : component cineraria_core_id_router_004
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                        --       src.ready
			src_valid          => id_router_006_src_valid,                                                        --          .valid
			src_data           => id_router_006_src_data,                                                         --          .data
			src_channel        => id_router_006_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                   --          .endofpacket
		);

	id_router_007 : component cineraria_core_id_router_004
		port map (
			sink_ready         => systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => systimer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                --       src.ready
			src_valid          => id_router_007_src_valid,                                                --          .valid
			src_data           => id_router_007_src_data,                                                 --          .data
			src_channel        => id_router_007_src_channel,                                              --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                           --          .endofpacket
		);

	id_router_008 : component cineraria_core_id_router_004
		port map (
			sink_ready         => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                           --       src.ready
			src_valid          => id_router_008_src_valid,                                           --          .valid
			src_data           => id_router_008_src_data,                                            --          .data
			src_channel        => id_router_008_src_channel,                                         --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                      --          .endofpacket
		);

	id_router_009 : component cineraria_core_id_router_004
		port map (
			sink_ready         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_7seg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                --       src.ready
			src_valid          => id_router_009_src_valid,                                                --          .valid
			src_data           => id_router_009_src_data,                                                 --          .data
			src_channel        => id_router_009_src_channel,                                              --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                           --          .endofpacket
		);

	id_router_010 : component cineraria_core_id_router_004
		port map (
			sink_ready         => psw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => psw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => psw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => psw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => psw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                           --       src.ready
			src_valid          => id_router_010_src_valid,                                           --          .valid
			src_data           => id_router_010_src_data,                                            --          .data
			src_channel        => id_router_010_src_channel,                                         --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                      --          .endofpacket
		);

	id_router_011 : component cineraria_core_id_router_004
		port map (
			sink_ready         => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dipsw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                             --       src.ready
			src_valid          => id_router_011_src_valid,                                             --          .valid
			src_data           => id_router_011_src_data,                                              --          .data
			src_channel        => id_router_011_src_channel,                                           --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                        --          .endofpacket
		);

	id_router_012 : component cineraria_core_id_router_004
		port map (
			sink_ready         => spu_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => spu_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => spu_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => spu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => spu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                           --       src.ready
			src_valid          => id_router_012_src_valid,                                           --          .valid
			src_data           => id_router_012_src_data,                                            --          .data
			src_channel        => id_router_012_src_channel,                                         --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                      --          .endofpacket
		);

	id_router_013 : component cineraria_core_id_router_004
		port map (
			sink_ready         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => mmcdma_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                              --       src.ready
			src_valid          => id_router_013_src_valid,                                              --          .valid
			src_data           => id_router_013_src_data,                                               --          .data
			src_channel        => id_router_013_src_channel,                                            --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                         --          .endofpacket
		);

	id_router_014 : component cineraria_core_id_router_004
		port map (
			sink_ready         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ps2_keyboard_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                                              --       src.ready
			src_valid          => id_router_014_src_valid,                                                              --          .valid
			src_data           => id_router_014_src_data,                                                               --          .data
			src_channel        => id_router_014_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                                         --          .endofpacket
		);

	id_router_015 : component cineraria_core_id_router_004
		port map (
			sink_ready         => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => gpio1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                             --       src.ready
			src_valid          => id_router_015_src_valid,                                             --          .valid
			src_data           => id_router_015_src_data,                                              --          .data
			src_channel        => id_router_015_src_channel,                                           --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                        --          .endofpacket
		);

	id_router_016 : component cineraria_core_id_router_004
		port map (
			sink_ready         => vga_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => vga_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => vga_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => vga_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                           --       src.ready
			src_valid          => id_router_016_src_valid,                                           --          .valid
			src_data           => id_router_016_src_data,                                            --          .data
			src_channel        => id_router_016_src_channel,                                         --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                      --          .endofpacket
		);

	id_router_017 : component cineraria_core_id_router_004
		port map (
			sink_ready         => blcon_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => blcon_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => blcon_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => blcon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => blcon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_40mhz_clk,                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_017_src_ready,                                             --       src.ready
			src_valid          => id_router_017_src_valid,                                             --          .valid
			src_data           => id_router_017_src_data,                                              --          .data
			src_channel        => id_router_017_src_channel,                                           --          .channel
			src_startofpacket  => id_router_017_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_017_src_endofpacket                                        --          .endofpacket
		);

	limiter : component cineraria_core_limiter
		generic map (
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			MAX_OUTSTANDING_RESPONSES => 9,
			PIPELINED                 => 0,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			VALID_WIDTH               => 4,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_100mhz_clk,                     --       clk.clk
			reset                  => rst_controller_001_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,              --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,              --          .valid
			cmd_sink_data          => addr_router_src_data,               --          .data
			cmd_sink_channel       => addr_router_src_channel,            --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,      --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,        --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,              --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,               --          .data
			cmd_src_channel        => limiter_cmd_src_channel,            --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,      --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,        --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,             --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,             --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,           --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,              --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket,     --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,       --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,              --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,              --          .valid
			rsp_src_data           => limiter_rsp_src_data,               --          .data
			rsp_src_channel        => limiter_rsp_src_channel,            --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,      --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,        --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data              -- cmd_valid.data
		);

	limiter_001 : component cineraria_core_limiter
		generic map (
			PKT_DEST_ID_H             => 104,
			PKT_DEST_ID_L             => 103,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			MAX_OUTSTANDING_RESPONSES => 10,
			PIPELINED                 => 0,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			VALID_WIDTH               => 4,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_100mhz_clk,                     --       clk.clk
			reset                  => rst_controller_001_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	limiter_002 : component cineraria_core_limiter_002
		generic map (
			PKT_DEST_ID_H             => 76,
			PKT_DEST_ID_L             => 73,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			MAX_OUTSTANDING_RESPONSES => 1,
			PIPELINED                 => 0,
			ST_DATA_W                 => 87,
			ST_CHANNEL_W              => 14,
			VALID_WIDTH               => 14,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 58,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_40mhz_clk,                      --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_004_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_004_src_valid,          --          .valid
			cmd_sink_data          => addr_router_004_src_data,           --          .data
			cmd_sink_channel       => addr_router_004_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_004_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_004_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_002_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_002_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_002_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_002_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_002_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_004_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_004_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_004_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_004_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_004_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_004_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_002_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_002_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_002_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_002_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_002_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_002_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_002_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component cineraria_core_burst_adapter
		generic map (
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 99,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			OUT_BYTE_CNT_H            => 76,
			OUT_BURSTWRAP_H           => 91,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 31,
			BURSTWRAP_CONST_VALUE     => 31
		)
		port map (
			clk                   => clk_100mhz_clk,                      --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,  -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_src_ready,              --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component cineraria_core_burst_adapter
		generic map (
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 99,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			OUT_BYTE_CNT_H            => 76,
			OUT_BURSTWRAP_H           => 91,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 31,
			BURSTWRAP_CONST_VALUE     => 31
		)
		port map (
			clk                   => clk_100mhz_clk,                          --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_001_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_001_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_001_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_001_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_001_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_001_src_ready,              --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	burst_adapter_002 : component cineraria_core_burst_adapter_002
		generic map (
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 81,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 76,
			PKT_BURST_SIZE_L          => 74,
			PKT_BURST_TYPE_H          => 78,
			PKT_BURST_TYPE_L          => 77,
			PKT_BURSTWRAP_H           => 73,
			PKT_BURSTWRAP_L           => 68,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 97,
			ST_CHANNEL_W              => 4,
			OUT_BYTE_CNT_H            => 57,
			OUT_BURSTWRAP_H           => 73,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 31,
			BURSTWRAP_CONST_VALUE     => 31
		)
		port map (
			clk                   => clk_100mhz_clk,                          --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_002_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_002_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_002_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_002_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_002_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_002_src_ready,              --          .ready
			source0_valid         => burst_adapter_002_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_002_source0_data,          --          .data
			source0_channel       => burst_adapter_002_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_002_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_002_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_002_source0_ready          --          .ready
		);

	burst_adapter_003 : component cineraria_core_burst_adapter
		generic map (
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 99,
			PKT_BYTE_CNT_H            => 85,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 94,
			PKT_BURST_SIZE_L          => 92,
			PKT_BURST_TYPE_H          => 96,
			PKT_BURST_TYPE_L          => 95,
			PKT_BURSTWRAP_H           => 91,
			PKT_BURSTWRAP_L           => 86,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 115,
			ST_CHANNEL_W              => 4,
			OUT_BYTE_CNT_H            => 76,
			OUT_BURSTWRAP_H           => 91,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 63,
			BURSTWRAP_CONST_VALUE     => 63
		)
		port map (
			clk                   => clk_100mhz_clk,                          --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_demux_001_src3_valid,           --     sink0.valid
			sink0_data            => cmd_xbar_demux_001_src3_data,            --          .data
			sink0_channel         => cmd_xbar_demux_001_src3_channel,         --          .channel
			sink0_startofpacket   => cmd_xbar_demux_001_src3_startofpacket,   --          .startofpacket
			sink0_endofpacket     => cmd_xbar_demux_001_src3_endofpacket,     --          .endofpacket
			sink0_ready           => cmd_xbar_demux_001_src3_ready,           --          .ready
			source0_valid         => burst_adapter_003_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_003_source0_data,          --          .data
			source0_channel       => burst_adapter_003_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_003_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_003_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_003_source0_ready          --          .ready
		);

	rst_controller : component cineraria_core_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk        => clk_40mhz_clk,                  --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component cineraria_core_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => sys_reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_100mhz_clk,                         --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_in1  => '0',                                    -- (terminated)
			reset_in2  => '0',                                    -- (terminated)
			reset_in3  => '0',                                    -- (terminated)
			reset_in4  => '0',                                    -- (terminated)
			reset_in5  => '0',                                    -- (terminated)
			reset_in6  => '0',                                    -- (terminated)
			reset_in7  => '0',                                    -- (terminated)
			reset_in8  => '0',                                    -- (terminated)
			reset_in9  => '0',                                    -- (terminated)
			reset_in10 => '0',                                    -- (terminated)
			reset_in11 => '0',                                    -- (terminated)
			reset_in12 => '0',                                    -- (terminated)
			reset_in13 => '0',                                    -- (terminated)
			reset_in14 => '0',                                    -- (terminated)
			reset_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component cineraria_core_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => sys_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_100mhz_clk,                     --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component cineraria_core_cmd_xbar_demux
		port map (
			clk                => clk_100mhz_clk,                     --        clk.clk
			reset              => rst_controller_001_reset_out_reset, --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,              --       sink.ready
			sink_channel       => limiter_cmd_src_channel,            --           .channel
			sink_data          => limiter_cmd_src_data,               --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,        --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,             -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,          --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,          --           .valid
			src0_data          => cmd_xbar_demux_src0_data,           --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,        --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket,  --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,    --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,          --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,          --           .valid
			src1_data          => cmd_xbar_demux_src1_data,           --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,        --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket,  --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,    --           .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,          --       src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,          --           .valid
			src2_data          => cmd_xbar_demux_src2_data,           --           .data
			src2_channel       => cmd_xbar_demux_src2_channel,        --           .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket,  --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket     --           .endofpacket
		);

	cmd_xbar_demux_001 : component cineraria_core_cmd_xbar_demux_001
		port map (
			clk                => clk_100mhz_clk,                        --        clk.clk
			reset              => rst_controller_001_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_001_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_001_cmd_src_channel,           --           .channel
			sink_data          => limiter_001_cmd_src_data,              --           .data
			sink_startofpacket => limiter_001_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_001_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_001_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --           .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --       src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --           .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --           .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --           .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_002 : component cineraria_core_cmd_xbar_demux_002
		port map (
			clk                => clk_100mhz_clk,                        --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_002_src_ready,             --      sink.ready
			sink_channel       => addr_router_002_src_channel,           --          .channel
			sink_data          => addr_router_002_src_data,              --          .data
			sink_startofpacket => addr_router_002_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_002_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_002_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_002_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_003 : component cineraria_core_cmd_xbar_demux_003
		port map (
			clk                => clk_100mhz_clk,                        --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_003_src_ready,             --      sink.ready
			sink_channel       => addr_router_003_src_channel,           --          .channel
			sink_data          => addr_router_003_src_data,              --          .data
			sink_startofpacket => addr_router_003_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_003_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_003_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_003_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component cineraria_core_cmd_xbar_mux
		port map (
			clk                 => clk_100mhz_clk,                        --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component cineraria_core_cmd_xbar_mux
		port map (
			clk                 => clk_100mhz_clk,                        --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component cineraria_core_cmd_xbar_mux_002
		port map (
			clk                 => clk_100mhz_clk,                        --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => width_adapter_src_ready,               --     sink0.ready
			sink0_valid         => width_adapter_src_valid,               --          .valid
			sink0_channel       => width_adapter_src_channel,             --          .channel
			sink0_data          => width_adapter_src_data,                --          .data
			sink0_startofpacket => width_adapter_src_startofpacket,       --          .startofpacket
			sink0_endofpacket   => width_adapter_src_endofpacket,         --          .endofpacket
			sink1_ready         => width_adapter_001_src_ready,           --     sink1.ready
			sink1_valid         => width_adapter_001_src_valid,           --          .valid
			sink1_channel       => width_adapter_001_src_channel,         --          .channel
			sink1_data          => width_adapter_001_src_data,            --          .data
			sink1_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink1_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink2_ready         => cmd_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => cmd_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => cmd_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => width_adapter_002_src_ready,           --     sink3.ready
			sink3_valid         => width_adapter_002_src_valid,           --          .valid
			sink3_channel       => width_adapter_002_src_channel,         --          .channel
			sink3_data          => width_adapter_002_src_data,            --          .data
			sink3_startofpacket => width_adapter_002_src_startofpacket,   --          .startofpacket
			sink3_endofpacket   => width_adapter_002_src_endofpacket      --          .endofpacket
		);

	rsp_xbar_demux : component cineraria_core_rsp_xbar_demux
		port map (
			clk                => clk_100mhz_clk,                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sink_ready         => id_router_src_ready,                --      sink.ready
			sink_channel       => id_router_src_channel,              --          .channel
			sink_data          => id_router_src_data,                 --          .data
			sink_startofpacket => id_router_src_startofpacket,        --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,          --          .endofpacket
			sink_valid(0)      => id_router_src_valid,                --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,          --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,          --          .valid
			src0_data          => rsp_xbar_demux_src0_data,           --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,          --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,          --          .valid
			src1_data          => rsp_xbar_demux_src1_data,           --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket     --          .endofpacket
		);

	rsp_xbar_demux_001 : component cineraria_core_rsp_xbar_demux
		port map (
			clk                => clk_100mhz_clk,                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component cineraria_core_rsp_xbar_demux_002
		port map (
			clk                => clk_100mhz_clk,                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_002_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_002_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_002_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_002_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_002_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_002_src2_endofpacket,   --          .endofpacket
			src3_ready         => rsp_xbar_demux_002_src3_ready,         --      src3.ready
			src3_valid         => rsp_xbar_demux_002_src3_valid,         --          .valid
			src3_data          => rsp_xbar_demux_002_src3_data,          --          .data
			src3_channel       => rsp_xbar_demux_002_src3_channel,       --          .channel
			src3_startofpacket => rsp_xbar_demux_002_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => rsp_xbar_demux_002_src3_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component cineraria_core_cmd_xbar_demux_003
		port map (
			clk                => clk_100mhz_clk,                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component cineraria_core_rsp_xbar_mux
		port map (
			clk                 => clk_100mhz_clk,                        --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => width_adapter_003_src_ready,           --     sink2.ready
			sink2_valid         => width_adapter_003_src_valid,           --          .valid
			sink2_channel       => width_adapter_003_src_channel,         --          .channel
			sink2_data          => width_adapter_003_src_data,            --          .data
			sink2_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink2_endofpacket   => width_adapter_003_src_endofpacket      --          .endofpacket
		);

	rsp_xbar_mux_001 : component cineraria_core_rsp_xbar_mux_001
		port map (
			clk                 => clk_100mhz_clk,                        --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => width_adapter_004_src_ready,           --     sink2.ready
			sink2_valid         => width_adapter_004_src_valid,           --          .valid
			sink2_channel       => width_adapter_004_src_channel,         --          .channel
			sink2_data          => width_adapter_004_src_data,            --          .data
			sink2_startofpacket => width_adapter_004_src_startofpacket,   --          .startofpacket
			sink2_endofpacket   => width_adapter_004_src_endofpacket,     --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_004 : component cineraria_core_cmd_xbar_demux_004
		port map (
			clk                 => clk_40mhz_clk,                          --        clk.clk
			reset               => rst_controller_reset_out_reset,         --  clk_reset.reset
			sink_ready          => limiter_002_cmd_src_ready,              --       sink.ready
			sink_channel        => limiter_002_cmd_src_channel,            --           .channel
			sink_data           => limiter_002_cmd_src_data,               --           .data
			sink_startofpacket  => limiter_002_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket    => limiter_002_cmd_src_endofpacket,        --           .endofpacket
			sink_valid          => limiter_002_cmd_valid_data,             -- sink_valid.data
			src0_ready          => cmd_xbar_demux_004_src0_ready,          --       src0.ready
			src0_valid          => cmd_xbar_demux_004_src0_valid,          --           .valid
			src0_data           => cmd_xbar_demux_004_src0_data,           --           .data
			src0_channel        => cmd_xbar_demux_004_src0_channel,        --           .channel
			src0_startofpacket  => cmd_xbar_demux_004_src0_startofpacket,  --           .startofpacket
			src0_endofpacket    => cmd_xbar_demux_004_src0_endofpacket,    --           .endofpacket
			src1_ready          => cmd_xbar_demux_004_src1_ready,          --       src1.ready
			src1_valid          => cmd_xbar_demux_004_src1_valid,          --           .valid
			src1_data           => cmd_xbar_demux_004_src1_data,           --           .data
			src1_channel        => cmd_xbar_demux_004_src1_channel,        --           .channel
			src1_startofpacket  => cmd_xbar_demux_004_src1_startofpacket,  --           .startofpacket
			src1_endofpacket    => cmd_xbar_demux_004_src1_endofpacket,    --           .endofpacket
			src2_ready          => cmd_xbar_demux_004_src2_ready,          --       src2.ready
			src2_valid          => cmd_xbar_demux_004_src2_valid,          --           .valid
			src2_data           => cmd_xbar_demux_004_src2_data,           --           .data
			src2_channel        => cmd_xbar_demux_004_src2_channel,        --           .channel
			src2_startofpacket  => cmd_xbar_demux_004_src2_startofpacket,  --           .startofpacket
			src2_endofpacket    => cmd_xbar_demux_004_src2_endofpacket,    --           .endofpacket
			src3_ready          => cmd_xbar_demux_004_src3_ready,          --       src3.ready
			src3_valid          => cmd_xbar_demux_004_src3_valid,          --           .valid
			src3_data           => cmd_xbar_demux_004_src3_data,           --           .data
			src3_channel        => cmd_xbar_demux_004_src3_channel,        --           .channel
			src3_startofpacket  => cmd_xbar_demux_004_src3_startofpacket,  --           .startofpacket
			src3_endofpacket    => cmd_xbar_demux_004_src3_endofpacket,    --           .endofpacket
			src4_ready          => cmd_xbar_demux_004_src4_ready,          --       src4.ready
			src4_valid          => cmd_xbar_demux_004_src4_valid,          --           .valid
			src4_data           => cmd_xbar_demux_004_src4_data,           --           .data
			src4_channel        => cmd_xbar_demux_004_src4_channel,        --           .channel
			src4_startofpacket  => cmd_xbar_demux_004_src4_startofpacket,  --           .startofpacket
			src4_endofpacket    => cmd_xbar_demux_004_src4_endofpacket,    --           .endofpacket
			src5_ready          => cmd_xbar_demux_004_src5_ready,          --       src5.ready
			src5_valid          => cmd_xbar_demux_004_src5_valid,          --           .valid
			src5_data           => cmd_xbar_demux_004_src5_data,           --           .data
			src5_channel        => cmd_xbar_demux_004_src5_channel,        --           .channel
			src5_startofpacket  => cmd_xbar_demux_004_src5_startofpacket,  --           .startofpacket
			src5_endofpacket    => cmd_xbar_demux_004_src5_endofpacket,    --           .endofpacket
			src6_ready          => cmd_xbar_demux_004_src6_ready,          --       src6.ready
			src6_valid          => cmd_xbar_demux_004_src6_valid,          --           .valid
			src6_data           => cmd_xbar_demux_004_src6_data,           --           .data
			src6_channel        => cmd_xbar_demux_004_src6_channel,        --           .channel
			src6_startofpacket  => cmd_xbar_demux_004_src6_startofpacket,  --           .startofpacket
			src6_endofpacket    => cmd_xbar_demux_004_src6_endofpacket,    --           .endofpacket
			src7_ready          => cmd_xbar_demux_004_src7_ready,          --       src7.ready
			src7_valid          => cmd_xbar_demux_004_src7_valid,          --           .valid
			src7_data           => cmd_xbar_demux_004_src7_data,           --           .data
			src7_channel        => cmd_xbar_demux_004_src7_channel,        --           .channel
			src7_startofpacket  => cmd_xbar_demux_004_src7_startofpacket,  --           .startofpacket
			src7_endofpacket    => cmd_xbar_demux_004_src7_endofpacket,    --           .endofpacket
			src8_ready          => cmd_xbar_demux_004_src8_ready,          --       src8.ready
			src8_valid          => cmd_xbar_demux_004_src8_valid,          --           .valid
			src8_data           => cmd_xbar_demux_004_src8_data,           --           .data
			src8_channel        => cmd_xbar_demux_004_src8_channel,        --           .channel
			src8_startofpacket  => cmd_xbar_demux_004_src8_startofpacket,  --           .startofpacket
			src8_endofpacket    => cmd_xbar_demux_004_src8_endofpacket,    --           .endofpacket
			src9_ready          => cmd_xbar_demux_004_src9_ready,          --       src9.ready
			src9_valid          => cmd_xbar_demux_004_src9_valid,          --           .valid
			src9_data           => cmd_xbar_demux_004_src9_data,           --           .data
			src9_channel        => cmd_xbar_demux_004_src9_channel,        --           .channel
			src9_startofpacket  => cmd_xbar_demux_004_src9_startofpacket,  --           .startofpacket
			src9_endofpacket    => cmd_xbar_demux_004_src9_endofpacket,    --           .endofpacket
			src10_ready         => cmd_xbar_demux_004_src10_ready,         --      src10.ready
			src10_valid         => cmd_xbar_demux_004_src10_valid,         --           .valid
			src10_data          => cmd_xbar_demux_004_src10_data,          --           .data
			src10_channel       => cmd_xbar_demux_004_src10_channel,       --           .channel
			src10_startofpacket => cmd_xbar_demux_004_src10_startofpacket, --           .startofpacket
			src10_endofpacket   => cmd_xbar_demux_004_src10_endofpacket,   --           .endofpacket
			src11_ready         => cmd_xbar_demux_004_src11_ready,         --      src11.ready
			src11_valid         => cmd_xbar_demux_004_src11_valid,         --           .valid
			src11_data          => cmd_xbar_demux_004_src11_data,          --           .data
			src11_channel       => cmd_xbar_demux_004_src11_channel,       --           .channel
			src11_startofpacket => cmd_xbar_demux_004_src11_startofpacket, --           .startofpacket
			src11_endofpacket   => cmd_xbar_demux_004_src11_endofpacket,   --           .endofpacket
			src12_ready         => cmd_xbar_demux_004_src12_ready,         --      src12.ready
			src12_valid         => cmd_xbar_demux_004_src12_valid,         --           .valid
			src12_data          => cmd_xbar_demux_004_src12_data,          --           .data
			src12_channel       => cmd_xbar_demux_004_src12_channel,       --           .channel
			src12_startofpacket => cmd_xbar_demux_004_src12_startofpacket, --           .startofpacket
			src12_endofpacket   => cmd_xbar_demux_004_src12_endofpacket,   --           .endofpacket
			src13_ready         => cmd_xbar_demux_004_src13_ready,         --      src13.ready
			src13_valid         => cmd_xbar_demux_004_src13_valid,         --           .valid
			src13_data          => cmd_xbar_demux_004_src13_data,          --           .data
			src13_channel       => cmd_xbar_demux_004_src13_channel,       --           .channel
			src13_startofpacket => cmd_xbar_demux_004_src13_startofpacket, --           .startofpacket
			src13_endofpacket   => cmd_xbar_demux_004_src13_endofpacket    --           .endofpacket
		);

	rsp_xbar_demux_004 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_017 : component cineraria_core_rsp_xbar_demux_004
		port map (
			clk                => clk_40mhz_clk,                         --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_017_src_ready,               --      sink.ready
			sink_channel       => id_router_017_src_channel,             --          .channel
			sink_data          => id_router_017_src_data,                --          .data
			sink_startofpacket => id_router_017_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_017_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_017_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_017_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_017_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_017_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_004 : component cineraria_core_rsp_xbar_mux_004
		port map (
			clk                  => clk_40mhz_clk,                         --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_004_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_004_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_004_src_data,             --          .data
			src_channel          => rsp_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_004_src0_ready,         --     sink0.ready
			sink0_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink0_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink0_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink0_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink1_ready          => rsp_xbar_demux_005_src0_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_006_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_007_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_008_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_009_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_010_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_010_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_011_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_011_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_012_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_012_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_013_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_013_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_014_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_015_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_016_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_016_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_017_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_017_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_017_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component cineraria_core_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 85,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 91,
			IN_PKT_BURSTWRAP_L            => 86,
			IN_PKT_BURST_SIZE_H           => 94,
			IN_PKT_BURST_SIZE_L           => 92,
			IN_PKT_RESPONSE_STATUS_H      => 114,
			IN_PKT_RESPONSE_STATUS_L      => 113,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 96,
			IN_PKT_BURST_TYPE_L           => 95,
			IN_ST_DATA_W                  => 115,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 67,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 76,
			OUT_PKT_BURST_SIZE_L          => 74,
			OUT_PKT_RESPONSE_STATUS_H     => 96,
			OUT_PKT_RESPONSE_STATUS_L     => 95,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 78,
			OUT_PKT_BURST_TYPE_L          => 77,
			OUT_ST_DATA_W                 => 97,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_100mhz_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset, -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src2_valid,          --      sink.valid
			in_channel           => cmd_xbar_demux_src2_channel,        --          .channel
			in_startofpacket     => cmd_xbar_demux_src2_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src2_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_demux_src2_ready,          --          .ready
			in_data              => cmd_xbar_demux_src2_data,           --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component cineraria_core_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 85,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 91,
			IN_PKT_BURSTWRAP_L            => 86,
			IN_PKT_BURST_SIZE_H           => 94,
			IN_PKT_BURST_SIZE_L           => 92,
			IN_PKT_RESPONSE_STATUS_H      => 114,
			IN_PKT_RESPONSE_STATUS_L      => 113,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 96,
			IN_PKT_BURST_TYPE_L           => 95,
			IN_ST_DATA_W                  => 115,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 67,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 76,
			OUT_PKT_BURST_SIZE_L          => 74,
			OUT_PKT_RESPONSE_STATUS_H     => 96,
			OUT_PKT_RESPONSE_STATUS_L     => 95,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 78,
			OUT_PKT_BURST_TYPE_L          => 77,
			OUT_ST_DATA_W                 => 97,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_100mhz_clk,                        --       clk.clk
			reset                => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src2_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src2_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src2_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src2_data,          --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_001_src_data,            --          .data
			out_channel          => width_adapter_001_src_channel,         --          .channel
			out_valid            => width_adapter_001_src_valid,           --          .valid
			out_ready            => width_adapter_001_src_ready,           --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_002 : component cineraria_core_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 85,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 91,
			IN_PKT_BURSTWRAP_L            => 86,
			IN_PKT_BURST_SIZE_H           => 94,
			IN_PKT_BURST_SIZE_L           => 92,
			IN_PKT_RESPONSE_STATUS_H      => 114,
			IN_PKT_RESPONSE_STATUS_L      => 113,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 96,
			IN_PKT_BURST_TYPE_L           => 95,
			IN_ST_DATA_W                  => 115,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 67,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 76,
			OUT_PKT_BURST_SIZE_L          => 74,
			OUT_PKT_RESPONSE_STATUS_H     => 96,
			OUT_PKT_RESPONSE_STATUS_L     => 95,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 78,
			OUT_PKT_BURST_TYPE_L          => 77,
			OUT_ST_DATA_W                 => 97,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_100mhz_clk,                        --       clk.clk
			reset                => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_003_src0_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_003_src0_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_003_src0_ready,         --          .ready
			in_data              => cmd_xbar_demux_003_src0_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_002_src_data,            --          .data
			out_channel          => width_adapter_002_src_channel,         --          .channel
			out_valid            => width_adapter_002_src_valid,           --          .valid
			out_ready            => width_adapter_002_src_ready,           --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_003 : component cineraria_core_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 67,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 73,
			IN_PKT_BURSTWRAP_L            => 68,
			IN_PKT_BURST_SIZE_H           => 76,
			IN_PKT_BURST_SIZE_L           => 74,
			IN_PKT_RESPONSE_STATUS_H      => 96,
			IN_PKT_RESPONSE_STATUS_L      => 95,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 78,
			IN_PKT_BURST_TYPE_L           => 77,
			IN_ST_DATA_W                  => 97,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 85,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 94,
			OUT_PKT_BURST_SIZE_L          => 92,
			OUT_PKT_RESPONSE_STATUS_H     => 114,
			OUT_PKT_RESPONSE_STATUS_L     => 113,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 96,
			OUT_PKT_BURST_TYPE_L          => 95,
			OUT_ST_DATA_W                 => 115,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_100mhz_clk,                        --       clk.clk
			reset                => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_002_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_002_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_002_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_002_src0_data,          --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_003_src_data,            --          .data
			out_channel          => width_adapter_003_src_channel,         --          .channel
			out_valid            => width_adapter_003_src_valid,           --          .valid
			out_ready            => width_adapter_003_src_ready,           --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_004 : component cineraria_core_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 67,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 73,
			IN_PKT_BURSTWRAP_L            => 68,
			IN_PKT_BURST_SIZE_H           => 76,
			IN_PKT_BURST_SIZE_L           => 74,
			IN_PKT_RESPONSE_STATUS_H      => 96,
			IN_PKT_RESPONSE_STATUS_L      => 95,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 78,
			IN_PKT_BURST_TYPE_L           => 77,
			IN_ST_DATA_W                  => 97,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 85,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 94,
			OUT_PKT_BURST_SIZE_L          => 92,
			OUT_PKT_RESPONSE_STATUS_H     => 114,
			OUT_PKT_RESPONSE_STATUS_L     => 113,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 96,
			OUT_PKT_BURST_TYPE_L          => 95,
			OUT_ST_DATA_W                 => 115,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_100mhz_clk,                        --       clk.clk
			reset                => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_002_src1_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_002_src1_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_002_src1_ready,         --          .ready
			in_data              => rsp_xbar_demux_002_src1_data,          --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_004_src_data,            --          .data
			out_channel          => width_adapter_004_src_channel,         --          .channel
			out_valid            => width_adapter_004_src_valid,           --          .valid
			out_ready            => width_adapter_004_src_ready,           --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_005 : component cineraria_core_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 67,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 73,
			IN_PKT_BURSTWRAP_L            => 68,
			IN_PKT_BURST_SIZE_H           => 76,
			IN_PKT_BURST_SIZE_L           => 74,
			IN_PKT_RESPONSE_STATUS_H      => 96,
			IN_PKT_RESPONSE_STATUS_L      => 95,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 78,
			IN_PKT_BURST_TYPE_L           => 77,
			IN_ST_DATA_W                  => 97,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 85,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 94,
			OUT_PKT_BURST_SIZE_L          => 92,
			OUT_PKT_RESPONSE_STATUS_H     => 114,
			OUT_PKT_RESPONSE_STATUS_L     => 113,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 96,
			OUT_PKT_BURST_TYPE_L          => 95,
			OUT_ST_DATA_W                 => 115,
			ST_CHANNEL_W                  => 4,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_100mhz_clk,                        --       clk.clk
			reset                => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			in_valid             => rsp_xbar_demux_002_src3_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_002_src3_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_002_src3_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_002_src3_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_002_src3_ready,         --          .ready
			in_data              => rsp_xbar_demux_002_src3_data,          --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_005_src_data,            --          .data
			out_channel          => width_adapter_005_src_channel,         --          .channel
			out_valid            => width_adapter_005_src_valid,           --          .valid
			out_ready            => width_adapter_005_src_ready,           --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	irq_mapper : component cineraria_core_irq_mapper
		port map (
			clk           => clk_100mhz_clk,                     --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,           -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,           -- receiver7.irq
			sender_irq    => nios2_fast_d_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver4_irq            --             sender.irq
		);

	irq_synchronizer_005 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_005_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver5_irq            --             sender.irq
		);

	irq_synchronizer_006 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_006_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver6_irq            --             sender.irq
		);

	irq_synchronizer_007 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_40mhz_clk,                      --       receiver_clk.clk
			sender_clk     => clk_100mhz_clk,                     --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_007_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver7_irq            --             sender.irq
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

	sdram_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_write;

	sdram_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_read;

	sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_byteenable;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	sysuart_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sysuart_s1_translator_avalon_anti_slave_0_write;

	sysuart_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sysuart_s1_translator_avalon_anti_slave_0_read;

	systimer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not systimer_s1_translator_avalon_anti_slave_0_write;

	led_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_s1_translator_avalon_anti_slave_0_write;

	led_7seg_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_7seg_s1_translator_avalon_anti_slave_0_write;

	psw_s1_translator_avalon_anti_slave_0_write_ports_inv <= not psw_s1_translator_avalon_anti_slave_0_write;

	gpio1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not gpio1_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of cineraria_core
