----------------------------------------------------------------------
-- TITLE : Loreley Compress Wave data Decoder
--
--     VERFASSER : S.OSAFUNE (J-7SYSTEM Works)
--     DATUM     : 2005/04/01 -> 2005/04/12 (HERSTELLUNG)
--               : 2005/04/12 (FESTSTELLUNG)
--
--               : 2006/01/05 �e�[�u����W��VHDL��
--               : 2006/09/24 �e�[�u�����g�p�I�v�V�����ǉ� (NEUBEARBEITUNG)
----------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity loreley_decoder is
	generic(
		CLOCK_EDGE		: std_logic := '1';	-- Rise edge drive clock
		RESET_LEVEL		: std_logic := '1';	-- Positive logic reset

		USE_DECODETABLE	: string := "ON";
		DECODE_TABLE	: string := "ROM_C352COMPRESS";
--		DECODE_TABLE	: string := "ROM_ALAWCOMPRESS";
--		DECODE_TABLE	: string := "ROM_ULAWCOMPRESS";
--		DECODE_TABLE	: string := "RAM";
		DEVICE_MAKER	: string := "ALTERA"
--		DEVICE_MAKER	: string := ""
	);
	port(
		clk				: in  std_logic;	-- system clock
		reset			: in  std_logic;	-- async reset

	--==== Decompresser I/F signal ===================================

		compress_data	: in  std_logic_vector(7 downto 0);
		decompress_data	: out std_logic_vector(15 downto 0);

	--==== System register I/F signal ================================

		dectable_rddata	: out std_logic_vector(31 downto 0);
		dectable_wrdata	: in  std_logic_vector(31 downto 0);
		dectable_write	: in  std_logic
	);
end loreley_decoder;

architecture RTL of loreley_decoder is
	type ROM_WORD is array(0 to 255) of std_logic_vector(15 downto 0);
	signal rom : ROM_WORD;
	signal compdata_reg		: std_logic_vector(7 downto 0);

	signal tableaddr_reg	: std_logic_vector(7 downto 0);
	signal tabledata_reg	: std_logic_vector(15 downto 0);
	signal tablewrite_sig	: std_logic;


	component loreley_simpledpram is
	generic(
		CLOCK_EDGE		: std_logic;
		RESET_LEVEL		: std_logic;
		ADDRESS_WIDTH	: integer;
		DATA_WIDTH		: integer;
		DEVICE_MAKER	: string
	);
	port(
		clk				: in  std_logic;
		reset			: in  std_logic :='0';

		rdaddress		: in  std_logic_vector(ADDRESS_WIDTH-1 downto 0);
		rddata			: out std_logic_vector(DATA_WIDTH-1 downto 0);
		wraddress		: in  std_logic_vector(ADDRESS_WIDTH-1 downto 0);
		wrdata			: in  std_logic_vector(DATA_WIDTH-1 downto 0);
		wrenable		: in  std_logic := '1'
	);
	end component;

begin

	-- �W�J�e�[�u����RAM�ŃC���X�^���X 
GEN_RAM : if (USE_DECODETABLE="ON" and DECODE_TABLE = "RAM") generate

	dectable_rddata(31 downto 24) <= (others=>'0');
	dectable_rddata(23 downto 16) <= tableaddr_reg;
	dectable_rddata(15 downto 0)  <= tabledata_reg;

	tablewrite_sig <= dectable_write and dectable_wrdata(24);

	process (clk,reset) begin
		if (reset=RESET_LEVEL) then
			tableaddr_reg <= (others=>'0');
			tabledata_reg <= (others=>'0');

		elsif (clk'event and clk=CLOCK_EDGE) then
			if (dectable_write='1') then
				tableaddr_reg <= dectable_wrdata(23 downto 16);
				tabledata_reg <= dectable_wrdata(15 downto 0);
			end if;

		end if;
	end process;

	U_ramtable : loreley_simpledpram
	generic map(
		CLOCK_EDGE		=> CLOCK_EDGE,
		RESET_LEVEL		=> RESET_LEVEL,
		ADDRESS_WIDTH	=> 8,
		DATA_WIDTH		=> 16,
		DEVICE_MAKER	=> DEVICE_MAKER
	)
	port map(
		clk			=> clk,
		reset		=> reset,

		rdaddress	=> compress_data,
		rddata		=> decompress_data,
		wraddress	=> dectable_wrdata(23 downto 16),
		wrdata		=> dectable_wrdata(15 downto 0),
		wrenable	=> tablewrite_sig
	);

	end generate;
GEN_TABLE : if (USE_DECODETABLE="ON" and DECODE_TABLE /= "RAM") generate

	dectable_rddata <= (others=>'X');

	process (clk) begin
		if (clk'event and clk=CLOCK_EDGE) then
			compdata_reg <= compress_data;
		end if;
	end process;

	decompress_data <= rom(CONV_INTEGER(compdata_reg));

	end generate;
GEN_UNUSE : if (USE_DECODETABLE /= "ON") generate

	dectable_rddata <= (others=>'X');
	decompress_data <= (others=>'X');

	end generate;


	-- C352 8bit�W�J�e�[�u�� 
GEN_ROM_C352 : if (DECODE_TABLE = "ROM_C352COMPRESS") generate

		rom(0  ) <= "0000000000000000";
		rom(1  ) <= "0000000000100000";
		rom(2  ) <= "0000000001000000";
		rom(3  ) <= "0000000001100000";
		rom(4  ) <= "0000000010000000";
		rom(5  ) <= "0000000010100000";
		rom(6  ) <= "0000000011000000";
		rom(7  ) <= "0000000011100000";
		rom(8  ) <= "0000000100000000";
		rom(9  ) <= "0000000100100000";
		rom(10 ) <= "0000000101000000";
		rom(11 ) <= "0000000101100000";
		rom(12 ) <= "0000000110000000";
		rom(13 ) <= "0000000110100000";
		rom(14 ) <= "0000000111000000";
		rom(15 ) <= "0000000111100000";
		rom(16 ) <= "0000001000100000";
		rom(17 ) <= "0000001001100000";
		rom(18 ) <= "0000001010100000";
		rom(19 ) <= "0000001011100000";
		rom(20 ) <= "0000001100100000";
		rom(21 ) <= "0000001101100000";
		rom(22 ) <= "0000001110100000";
		rom(23 ) <= "0000001111100000";
		rom(24 ) <= "0000010001100001";
		rom(25 ) <= "0000010011100001";
		rom(26 ) <= "0000010101100001";
		rom(27 ) <= "0000010111100001";
		rom(28 ) <= "0000011001100001";
		rom(29 ) <= "0000011011100001";
		rom(30 ) <= "0000011101100001";
		rom(31 ) <= "0000011111100001";
		rom(32 ) <= "0000100001100010";
		rom(33 ) <= "0000100011100010";
		rom(34 ) <= "0000100101100010";
		rom(35 ) <= "0000100111100010";
		rom(36 ) <= "0000101001100010";
		rom(37 ) <= "0000101011100010";
		rom(38 ) <= "0000101101100010";
		rom(39 ) <= "0000101111100010";
		rom(40 ) <= "0000110001100011";
		rom(41 ) <= "0000110011100011";
		rom(42 ) <= "0000110101100011";
		rom(43 ) <= "0000110111100011";
		rom(44 ) <= "0000111001100011";
		rom(45 ) <= "0000111011100011";
		rom(46 ) <= "0000111101100011";
		rom(47 ) <= "0000111111100011";
		rom(48 ) <= "0001000011100100";
		rom(49 ) <= "0001000111100100";
		rom(50 ) <= "0001001011100100";
		rom(51 ) <= "0001001111100100";
		rom(52 ) <= "0001010011100101";
		rom(53 ) <= "0001010111100101";
		rom(54 ) <= "0001011011100101";
		rom(55 ) <= "0001011111100101";
		rom(56 ) <= "0001100011100110";
		rom(57 ) <= "0001100111100110";
		rom(58 ) <= "0001101011100110";
		rom(59 ) <= "0001101111100110";
		rom(60 ) <= "0001110011100111";
		rom(61 ) <= "0001110111100111";
		rom(62 ) <= "0001111011100111";
		rom(63 ) <= "0001111111100111";
		rom(64 ) <= "0010000011101000";
		rom(65 ) <= "0010000111101000";
		rom(66 ) <= "0010001011101000";
		rom(67 ) <= "0010001111101000";
		rom(68 ) <= "0010010011101001";
		rom(69 ) <= "0010010111101001";
		rom(70 ) <= "0010011011101001";
		rom(71 ) <= "0010011111101001";
		rom(72 ) <= "0010100011101010";
		rom(73 ) <= "0010100111101010";
		rom(74 ) <= "0010101011101010";
		rom(75 ) <= "0010101111101010";
		rom(76 ) <= "0010110011101011";
		rom(77 ) <= "0010110111101011";
		rom(78 ) <= "0010111011101011";
		rom(79 ) <= "0010111111101011";
		rom(80 ) <= "0011000011101100";
		rom(81 ) <= "0011000111101100";
		rom(82 ) <= "0011001011101100";
		rom(83 ) <= "0011001111101100";
		rom(84 ) <= "0011010011101101";
		rom(85 ) <= "0011010111101101";
		rom(86 ) <= "0011011011101101";
		rom(87 ) <= "0011011111101101";
		rom(88 ) <= "0011100011101110";
		rom(89 ) <= "0011100111101110";
		rom(90 ) <= "0011101011101110";
		rom(91 ) <= "0011101111101110";
		rom(92 ) <= "0011110011101111";
		rom(93 ) <= "0011110111101111";
		rom(94 ) <= "0011111011101111";
		rom(95 ) <= "0011111111101111";
		rom(96 ) <= "0100000011110000";
		rom(97 ) <= "0100000111110000";
		rom(98 ) <= "0100001011110000";
		rom(99 ) <= "0100001111110000";
		rom(100) <= "0100010111110001";
		rom(101) <= "0100011111110001";
		rom(102) <= "0100100111110010";
		rom(103) <= "0100101111110010";
		rom(104) <= "0100110111110011";
		rom(105) <= "0100111111110011";
		rom(106) <= "0101000111110100";
		rom(107) <= "0101001111110100";
		rom(108) <= "0101010111110101";
		rom(109) <= "0101011111110101";
		rom(110) <= "0101100111110110";
		rom(111) <= "0101101111110110";
		rom(112) <= "0101110111110111";
		rom(113) <= "0101111111110111";
		rom(114) <= "0110000111111000";
		rom(115) <= "0110001111111000";
		rom(116) <= "0110010111111001";
		rom(117) <= "0110011111111001";
		rom(118) <= "0110100111111010";
		rom(119) <= "0110101111111010";
		rom(120) <= "0110110111111011";
		rom(121) <= "0110111111111011";
		rom(122) <= "0111000111111100";
		rom(123) <= "0111001111111100";
		rom(124) <= "0111010111111101";
		rom(125) <= "0111011111111101";
		rom(126) <= "0111100111111110";
		rom(127) <= "0111111111111111";
		rom(128) <= "1000000000000000";
		rom(129) <= "1000011000000001";
		rom(130) <= "1000100000000010";
		rom(131) <= "1000101000000010";
		rom(132) <= "1000110000000011";
		rom(133) <= "1000111000000011";
		rom(134) <= "1001000000000100";
		rom(135) <= "1001001000000100";
		rom(136) <= "1001010000000101";
		rom(137) <= "1001011000000101";
		rom(138) <= "1001100000000110";
		rom(139) <= "1001101000000110";
		rom(140) <= "1001110000000111";
		rom(141) <= "1001111000000111";
		rom(142) <= "1010000000001000";
		rom(143) <= "1010001000001000";
		rom(144) <= "1010010000001001";
		rom(145) <= "1010011000001001";
		rom(146) <= "1010100000001010";
		rom(147) <= "1010101000001010";
		rom(148) <= "1010110000001011";
		rom(149) <= "1010111000001011";
		rom(150) <= "1011000000001100";
		rom(151) <= "1011001000001100";
		rom(152) <= "1011010000001101";
		rom(153) <= "1011011000001101";
		rom(154) <= "1011100000101110";
		rom(155) <= "1011101000001110";
		rom(156) <= "1011110000001111";
		rom(157) <= "1011110100001111";
		rom(158) <= "1011111000001111";
		rom(159) <= "1011111100001111";
		rom(160) <= "1100000000010000";
		rom(161) <= "1100000100010000";
		rom(162) <= "1100001000010000";
		rom(163) <= "1100001100010000";
		rom(164) <= "1100010000010001";
		rom(165) <= "1100010100010001";
		rom(166) <= "1100011000010001";
		rom(167) <= "1100011100010001";
		rom(168) <= "1100100000010010";
		rom(169) <= "1100100100010010";
		rom(170) <= "1100101000010010";
		rom(171) <= "1100101100010010";
		rom(172) <= "1100110000010011";
		rom(173) <= "1100110100010011";
		rom(174) <= "1100111000010011";
		rom(175) <= "1100111100010011";
		rom(176) <= "1101000000010100";
		rom(177) <= "1101000100010100";
		rom(178) <= "1101001000010100";
		rom(179) <= "1101001100010100";
		rom(180) <= "1101010000010101";
		rom(181) <= "1101010100010101";
		rom(182) <= "1101011000010101";
		rom(183) <= "1101011100010101";
		rom(184) <= "1101100000010110";
		rom(185) <= "1101100100010110";
		rom(186) <= "1101101000010110";
		rom(187) <= "1101101100010110";
		rom(188) <= "1101110000010111";
		rom(189) <= "1101110100010111";
		rom(190) <= "1101111000010111";
		rom(191) <= "1101111100010111";
		rom(192) <= "1110000000011000";
		rom(193) <= "1110000100011000";
		rom(194) <= "1110001000011000";
		rom(195) <= "1110001100011000";
		rom(196) <= "1110010000011001";
		rom(197) <= "1110010100011001";
		rom(198) <= "1110011000011001";
		rom(199) <= "1110011100011001";
		rom(200) <= "1110100000011010";
		rom(201) <= "1110100100011010";
		rom(202) <= "1110101000011010";
		rom(203) <= "1110101100011010";
		rom(204) <= "1110110000011011";
		rom(205) <= "1110110100011011";
		rom(206) <= "1110111000011011";
		rom(207) <= "1110111100011011";
		rom(208) <= "1111000000011100";
		rom(209) <= "1111000010011100";
		rom(210) <= "1111000100011100";
		rom(211) <= "1111000110011100";
		rom(212) <= "1111001000011100";
		rom(213) <= "1111001010011100";
		rom(214) <= "1111001100011100";
		rom(215) <= "1111001110011100";
		rom(216) <= "1111010000011101";
		rom(217) <= "1111010010011101";
		rom(218) <= "1111010100011101";
		rom(219) <= "1111010110011101";
		rom(220) <= "1111011000011101";
		rom(221) <= "1111011010011101";
		rom(222) <= "1111011100011101";
		rom(223) <= "1111011110011101";
		rom(224) <= "1111100000011110";
		rom(225) <= "1111100010011110";
		rom(226) <= "1111100100011110";
		rom(227) <= "1111100110011110";
		rom(228) <= "1111101000011110";
		rom(229) <= "1111101010011110";
		rom(230) <= "1111101100011110";
		rom(231) <= "1111101110011110";
		rom(232) <= "1111110000011111";
		rom(233) <= "1111110001011111";
		rom(234) <= "1111110010011111";
		rom(235) <= "1111110011011111";
		rom(236) <= "1111110100011111";
		rom(237) <= "1111110101011111";
		rom(238) <= "1111110110011111";
		rom(239) <= "1111110111011111";
		rom(240) <= "1111111000011111";
		rom(241) <= "1111111000111111";
		rom(242) <= "1111111001011111";
		rom(243) <= "1111111001111111";
		rom(244) <= "1111111010011111";
		rom(245) <= "1111111010111111";
		rom(246) <= "1111111011011111";
		rom(247) <= "1111111011111111";
		rom(248) <= "1111111100011111";
		rom(249) <= "1111111100111111";
		rom(250) <= "1111111101011111";
		rom(251) <= "1111111101111111";
		rom(252) <= "1111111110011111";
		rom(253) <= "1111111110111111";
		rom(254) <= "1111111111011111";
		rom(255) <= "1111111111111111";

	end generate;


	-- A-law 8bit�W�J�e�[�u�� 
GEN_ROM_ALAW : if (DECODE_TABLE = "ROM_ALAWCOMPRESS") generate

		rom(0  ) <= "1110101010000000";
		rom(1  ) <= "1110101110000000";
		rom(2  ) <= "1110100010000000";
		rom(3  ) <= "1110100110000000";
		rom(4  ) <= "1110111010000000";
		rom(5  ) <= "1110111110000000";
		rom(6  ) <= "1110110010000000";
		rom(7  ) <= "1110110110000000";
		rom(8  ) <= "1110001010000000";
		rom(9  ) <= "1110001110000000";
		rom(10 ) <= "1110000010000000";
		rom(11 ) <= "1110000110000000";
		rom(12 ) <= "1110011010000000";
		rom(13 ) <= "1110011110000000";
		rom(14 ) <= "1110010010000000";
		rom(15 ) <= "1110010110000000";
		rom(16 ) <= "1111010101000000";
		rom(17 ) <= "1111010111000000";
		rom(18 ) <= "1111010001000000";
		rom(19 ) <= "1111010011000000";
		rom(20 ) <= "1111011101000000";
		rom(21 ) <= "1111011111000000";
		rom(22 ) <= "1111011001000000";
		rom(23 ) <= "1111011011000000";
		rom(24 ) <= "1111000101000000";
		rom(25 ) <= "1111000111000000";
		rom(26 ) <= "1111000001000000";
		rom(27 ) <= "1111000011000000";
		rom(28 ) <= "1111001101000000";
		rom(29 ) <= "1111001111000000";
		rom(30 ) <= "1111001001000000";
		rom(31 ) <= "1111001011000000";
		rom(32 ) <= "1010101000000000";
		rom(33 ) <= "1010111000000000";
		rom(34 ) <= "1010001000000000";
		rom(35 ) <= "1010011000000000";
		rom(36 ) <= "1011101000000000";
		rom(37 ) <= "1011111000000000";
		rom(38 ) <= "1011001000000000";
		rom(39 ) <= "1011011000000000";
		rom(40 ) <= "1000101000000000";
		rom(41 ) <= "1000111000000000";
		rom(42 ) <= "1000001000000000";
		rom(43 ) <= "1000011000000000";
		rom(44 ) <= "1001101000000000";
		rom(45 ) <= "1001111000000000";
		rom(46 ) <= "1001001000000000";
		rom(47 ) <= "1001011000000000";
		rom(48 ) <= "1101010100000000";
		rom(49 ) <= "1101011100000000";
		rom(50 ) <= "1101000100000000";
		rom(51 ) <= "1101001100000000";
		rom(52 ) <= "1101110100000000";
		rom(53 ) <= "1101111100000000";
		rom(54 ) <= "1101100100000000";
		rom(55 ) <= "1101101100000000";
		rom(56 ) <= "1100010100000000";
		rom(57 ) <= "1100011100000000";
		rom(58 ) <= "1100000100000000";
		rom(59 ) <= "1100001100000000";
		rom(60 ) <= "1100110100000000";
		rom(61 ) <= "1100111100000000";
		rom(62 ) <= "1100100100000000";
		rom(63 ) <= "1100101100000000";
		rom(64 ) <= "1111111010101000";
		rom(65 ) <= "1111111010111000";
		rom(66 ) <= "1111111010001000";
		rom(67 ) <= "1111111010011000";
		rom(68 ) <= "1111111011101000";
		rom(69 ) <= "1111111011111000";
		rom(70 ) <= "1111111011001000";
		rom(71 ) <= "1111111011011000";
		rom(72 ) <= "1111111000101000";
		rom(73 ) <= "1111111000111000";
		rom(74 ) <= "1111111000001000";
		rom(75 ) <= "1111111000011000";
		rom(76 ) <= "1111111001101000";
		rom(77 ) <= "1111111001111000";
		rom(78 ) <= "1111111001001000";
		rom(79 ) <= "1111111001011000";
		rom(80 ) <= "1111111110101000";
		rom(81 ) <= "1111111110111000";
		rom(82 ) <= "1111111110001000";
		rom(83 ) <= "1111111110011000";
		rom(84 ) <= "1111111111101000";
		rom(85 ) <= "1111111111111000";
		rom(86 ) <= "1111111111001000";
		rom(87 ) <= "1111111111011000";
		rom(88 ) <= "1111111100101000";
		rom(89 ) <= "1111111100111000";
		rom(90 ) <= "1111111100001000";
		rom(91 ) <= "1111111100011000";
		rom(92 ) <= "1111111101101000";
		rom(93 ) <= "1111111101111000";
		rom(94 ) <= "1111111101001000";
		rom(95 ) <= "1111111101011000";
		rom(96 ) <= "1111101010100000";
		rom(97 ) <= "1111101011100000";
		rom(98 ) <= "1111101000100000";
		rom(99 ) <= "1111101001100000";
		rom(100) <= "1111101110100000";
		rom(101) <= "1111101111100000";
		rom(102) <= "1111101100100000";
		rom(103) <= "1111101101100000";
		rom(104) <= "1111100010100000";
		rom(105) <= "1111100011100000";
		rom(106) <= "1111100000100000";
		rom(107) <= "1111100001100000";
		rom(108) <= "1111100110100000";
		rom(109) <= "1111100111100000";
		rom(110) <= "1111100100100000";
		rom(111) <= "1111100101100000";
		rom(112) <= "1111110101010000";
		rom(113) <= "1111110101110000";
		rom(114) <= "1111110100010000";
		rom(115) <= "1111110100110000";
		rom(116) <= "1111110111010000";
		rom(117) <= "1111110111110000";
		rom(118) <= "1111110110010000";
		rom(119) <= "1111110110110000";
		rom(120) <= "1111110001010000";
		rom(121) <= "1111110001110000";
		rom(122) <= "1111110000010000";
		rom(123) <= "1111110000110000";
		rom(124) <= "1111110011010000";
		rom(125) <= "1111110011110000";
		rom(126) <= "1111110010010000";
		rom(127) <= "1111110010110000";
		rom(128) <= "0001010110000000";
		rom(129) <= "0001010010000000";
		rom(130) <= "0001011110000000";
		rom(131) <= "0001011010000000";
		rom(132) <= "0001000110000000";
		rom(133) <= "0001000010000000";
		rom(134) <= "0001001110000000";
		rom(135) <= "0001001010000000";
		rom(136) <= "0001110110000000";
		rom(137) <= "0001110010000000";
		rom(138) <= "0001111110000000";
		rom(139) <= "0001111010000000";
		rom(140) <= "0001100110000000";
		rom(141) <= "0001100010000000";
		rom(142) <= "0001101110000000";
		rom(143) <= "0001101010000000";
		rom(144) <= "0000101011000000";
		rom(145) <= "0000101001000000";
		rom(146) <= "0000101111000000";
		rom(147) <= "0000101101000000";
		rom(148) <= "0000100011000000";
		rom(149) <= "0000100001000000";
		rom(150) <= "0000100111000000";
		rom(151) <= "0000100101000000";
		rom(152) <= "0000111011000000";
		rom(153) <= "0000111001000000";
		rom(154) <= "0000111111000000";
		rom(155) <= "0000111101000000";
		rom(156) <= "0000110011000000";
		rom(157) <= "0000110001000000";
		rom(158) <= "0000110111000000";
		rom(159) <= "0000110101000000";
		rom(160) <= "0101011000000000";
		rom(161) <= "0101001000000000";
		rom(162) <= "0101111000000000";
		rom(163) <= "0101101000000000";
		rom(164) <= "0100011000000000";
		rom(165) <= "0100001000000000";
		rom(166) <= "0100111000000000";
		rom(167) <= "0100101000000000";
		rom(168) <= "0111011000000000";
		rom(169) <= "0111001000000000";
		rom(170) <= "0111111000000000";
		rom(171) <= "0111101000000000";
		rom(172) <= "0110011000000000";
		rom(173) <= "0110001000000000";
		rom(174) <= "0110111000000000";
		rom(175) <= "0110101000000000";
		rom(176) <= "0010101100000000";
		rom(177) <= "0010100100000000";
		rom(178) <= "0010111100000000";
		rom(179) <= "0010110100000000";
		rom(180) <= "0010001100000000";
		rom(181) <= "0010000100000000";
		rom(182) <= "0010011100000000";
		rom(183) <= "0010010100000000";
		rom(184) <= "0011101100000000";
		rom(185) <= "0011100100000000";
		rom(186) <= "0011111100000000";
		rom(187) <= "0011110100000000";
		rom(188) <= "0011001100000000";
		rom(189) <= "0011000100000000";
		rom(190) <= "0011011100000000";
		rom(191) <= "0011010100000000";
		rom(192) <= "0000000101011000";
		rom(193) <= "0000000101001000";
		rom(194) <= "0000000101111000";
		rom(195) <= "0000000101101000";
		rom(196) <= "0000000100011000";
		rom(197) <= "0000000100001000";
		rom(198) <= "0000000100111000";
		rom(199) <= "0000000100101000";
		rom(200) <= "0000000111011000";
		rom(201) <= "0000000111001000";
		rom(202) <= "0000000111111000";
		rom(203) <= "0000000111101000";
		rom(204) <= "0000000110011000";
		rom(205) <= "0000000110001000";
		rom(206) <= "0000000110111000";
		rom(207) <= "0000000110101000";
		rom(208) <= "0000000001011000";
		rom(209) <= "0000000001001000";
		rom(210) <= "0000000001111000";
		rom(211) <= "0000000001101000";
		rom(212) <= "0000000000011000";
		rom(213) <= "0000000000001000";
		rom(214) <= "0000000000111000";
		rom(215) <= "0000000000101000";
		rom(216) <= "0000000011011000";
		rom(217) <= "0000000011001000";
		rom(218) <= "0000000011111000";
		rom(219) <= "0000000011101000";
		rom(220) <= "0000000010011000";
		rom(221) <= "0000000010001000";
		rom(222) <= "0000000010111000";
		rom(223) <= "0000000010101000";
		rom(224) <= "0000010101100000";
		rom(225) <= "0000010100100000";
		rom(226) <= "0000010111100000";
		rom(227) <= "0000010110100000";
		rom(228) <= "0000010001100000";
		rom(229) <= "0000010000100000";
		rom(230) <= "0000010011100000";
		rom(231) <= "0000010010100000";
		rom(232) <= "0000011101100000";
		rom(233) <= "0000011100100000";
		rom(234) <= "0000011111100000";
		rom(235) <= "0000011110100000";
		rom(236) <= "0000011001100000";
		rom(237) <= "0000011000100000";
		rom(238) <= "0000011011100000";
		rom(239) <= "0000011010100000";
		rom(240) <= "0000001010110000";
		rom(241) <= "0000001010010000";
		rom(242) <= "0000001011110000";
		rom(243) <= "0000001011010000";
		rom(244) <= "0000001000110000";
		rom(245) <= "0000001000010000";
		rom(246) <= "0000001001110000";
		rom(247) <= "0000001001010000";
		rom(248) <= "0000001110110000";
		rom(249) <= "0000001110010000";
		rom(250) <= "0000001111110000";
		rom(251) <= "0000001111010000";
		rom(252) <= "0000001100110000";
		rom(253) <= "0000001100010000";
		rom(254) <= "0000001101110000";
		rom(255) <= "0000001101010000";

	end generate;


	-- ��-law 8bit�W�J�e�[�u�� 
GEN_ROM_ULAW : if (DECODE_TABLE = "ROM_ULAWCOMPRESS") generate

		rom(0  ) <= "1000001010000100";
		rom(1  ) <= "1000011010000100";
		rom(2  ) <= "1000101010000100";
		rom(3  ) <= "1000111010000100";
		rom(4  ) <= "1001001010000100";
		rom(5  ) <= "1001011010000100";
		rom(6  ) <= "1001101010000100";
		rom(7  ) <= "1001111010000100";
		rom(8  ) <= "1010001010000100";
		rom(9  ) <= "1010011010000100";
		rom(10 ) <= "1010101010000100";
		rom(11 ) <= "1010111010000100";
		rom(12 ) <= "1011001010000100";
		rom(13 ) <= "1011011010000100";
		rom(14 ) <= "1011101010000100";
		rom(15 ) <= "1011111010000100";
		rom(16 ) <= "1100000110000100";
		rom(17 ) <= "1100001110000100";
		rom(18 ) <= "1100010110000100";
		rom(19 ) <= "1100011110000100";
		rom(20 ) <= "1100100110000100";
		rom(21 ) <= "1100101110000100";
		rom(22 ) <= "1100110110000100";
		rom(23 ) <= "1100111110000100";
		rom(24 ) <= "1101000110000100";
		rom(25 ) <= "1101001110000100";
		rom(26 ) <= "1101010110000100";
		rom(27 ) <= "1101011110000100";
		rom(28 ) <= "1101100110000100";
		rom(29 ) <= "1101101110000100";
		rom(30 ) <= "1101110110000100";
		rom(31 ) <= "1101111110000100";
		rom(32 ) <= "1110000100000100";
		rom(33 ) <= "1110001000000100";
		rom(34 ) <= "1110001100000100";
		rom(35 ) <= "1110010000000100";
		rom(36 ) <= "1110010100000100";
		rom(37 ) <= "1110011000000100";
		rom(38 ) <= "1110011100000100";
		rom(39 ) <= "1110100000000100";
		rom(40 ) <= "1110100100000100";
		rom(41 ) <= "1110101000000100";
		rom(42 ) <= "1110101100000100";
		rom(43 ) <= "1110110000000100";
		rom(44 ) <= "1110110100000100";
		rom(45 ) <= "1110111000000100";
		rom(46 ) <= "1110111100000100";
		rom(47 ) <= "1111000000000100";
		rom(48 ) <= "1111000011000100";
		rom(49 ) <= "1111000101000100";
		rom(50 ) <= "1111000111000100";
		rom(51 ) <= "1111001001000100";
		rom(52 ) <= "1111001011000100";
		rom(53 ) <= "1111001101000100";
		rom(54 ) <= "1111001111000100";
		rom(55 ) <= "1111010001000100";
		rom(56 ) <= "1111010011000100";
		rom(57 ) <= "1111010101000100";
		rom(58 ) <= "1111010111000100";
		rom(59 ) <= "1111011001000100";
		rom(60 ) <= "1111011011000100";
		rom(61 ) <= "1111011101000100";
		rom(62 ) <= "1111011111000100";
		rom(63 ) <= "1111100001000100";
		rom(64 ) <= "1111100010100100";
		rom(65 ) <= "1111100011100100";
		rom(66 ) <= "1111100100100100";
		rom(67 ) <= "1111100101100100";
		rom(68 ) <= "1111100110100100";
		rom(69 ) <= "1111100111100100";
		rom(70 ) <= "1111101000100100";
		rom(71 ) <= "1111101001100100";
		rom(72 ) <= "1111101010100100";
		rom(73 ) <= "1111101011100100";
		rom(74 ) <= "1111101100100100";
		rom(75 ) <= "1111101101100100";
		rom(76 ) <= "1111101110100100";
		rom(77 ) <= "1111101111100100";
		rom(78 ) <= "1111110000100100";
		rom(79 ) <= "1111110001100100";
		rom(80 ) <= "1111110010010100";
		rom(81 ) <= "1111110010110100";
		rom(82 ) <= "1111110011010100";
		rom(83 ) <= "1111110011110100";
		rom(84 ) <= "1111110100010100";
		rom(85 ) <= "1111110100110100";
		rom(86 ) <= "1111110101010100";
		rom(87 ) <= "1111110101110100";
		rom(88 ) <= "1111110110010100";
		rom(89 ) <= "1111110110110100";
		rom(90 ) <= "1111110111010100";
		rom(91 ) <= "1111110111110100";
		rom(92 ) <= "1111111000010100";
		rom(93 ) <= "1111111000110100";
		rom(94 ) <= "1111111001010100";
		rom(95 ) <= "1111111001110100";
		rom(96 ) <= "1111111010001100";
		rom(97 ) <= "1111111010011100";
		rom(98 ) <= "1111111010101100";
		rom(99 ) <= "1111111010111100";
		rom(100) <= "1111111011001100";
		rom(101) <= "1111111011011100";
		rom(102) <= "1111111011101100";
		rom(103) <= "1111111011111100";
		rom(104) <= "1111111100001100";
		rom(105) <= "1111111100011100";
		rom(106) <= "1111111100101100";
		rom(107) <= "1111111100111100";
		rom(108) <= "1111111101001100";
		rom(109) <= "1111111101011100";
		rom(110) <= "1111111101101100";
		rom(111) <= "1111111101111100";
		rom(112) <= "1111111110001000";
		rom(113) <= "1111111110010000";
		rom(114) <= "1111111110011000";
		rom(115) <= "1111111110100000";
		rom(116) <= "1111111110101000";
		rom(117) <= "1111111110110000";
		rom(118) <= "1111111110111000";
		rom(119) <= "1111111111000000";
		rom(120) <= "1111111111001000";
		rom(121) <= "1111111111010000";
		rom(122) <= "1111111111011000";
		rom(123) <= "1111111111100000";
		rom(124) <= "1111111111101000";
		rom(125) <= "1111111111110000";
		rom(126) <= "1111111111111000";
		rom(127) <= "0000000000000000";
		rom(128) <= "0111110101111100";
		rom(129) <= "0111100101111100";
		rom(130) <= "0111010101111100";
		rom(131) <= "0111000101111100";
		rom(132) <= "0110110101111100";
		rom(133) <= "0110100101111100";
		rom(134) <= "0110010101111100";
		rom(135) <= "0110000101111100";
		rom(136) <= "0101110101111100";
		rom(137) <= "0101100101111100";
		rom(138) <= "0101010101111100";
		rom(139) <= "0101000101111100";
		rom(140) <= "0100110101111100";
		rom(141) <= "0100100101111100";
		rom(142) <= "0100010101111100";
		rom(143) <= "0100000101111100";
		rom(144) <= "0011111001111100";
		rom(145) <= "0011110001111100";
		rom(146) <= "0011101001111100";
		rom(147) <= "0011100001111100";
		rom(148) <= "0011011001111100";
		rom(149) <= "0011010001111100";
		rom(150) <= "0011001001111100";
		rom(151) <= "0011000001111100";
		rom(152) <= "0010111001111100";
		rom(153) <= "0010110001111100";
		rom(154) <= "0010101001111100";
		rom(155) <= "0010100001111100";
		rom(156) <= "0010011001111100";
		rom(157) <= "0010010001111100";
		rom(158) <= "0010001001111100";
		rom(159) <= "0010000001111100";
		rom(160) <= "0001111011111100";
		rom(161) <= "0001110111111100";
		rom(162) <= "0001110011111100";
		rom(163) <= "0001101111111100";
		rom(164) <= "0001101011111100";
		rom(165) <= "0001100111111100";
		rom(166) <= "0001100011111100";
		rom(167) <= "0001011111111100";
		rom(168) <= "0001011011111100";
		rom(169) <= "0001010111111100";
		rom(170) <= "0001010011111100";
		rom(171) <= "0001001111111100";
		rom(172) <= "0001001011111100";
		rom(173) <= "0001000111111100";
		rom(174) <= "0001000011111100";
		rom(175) <= "0000111111111100";
		rom(176) <= "0000111100111100";
		rom(177) <= "0000111010111100";
		rom(178) <= "0000111000111100";
		rom(179) <= "0000110110111100";
		rom(180) <= "0000110100111100";
		rom(181) <= "0000110010111100";
		rom(182) <= "0000110000111100";
		rom(183) <= "0000101110111100";
		rom(184) <= "0000101100111100";
		rom(185) <= "0000101010111100";
		rom(186) <= "0000101000111100";
		rom(187) <= "0000100110111100";
		rom(188) <= "0000100100111100";
		rom(189) <= "0000100010111100";
		rom(190) <= "0000100000111100";
		rom(191) <= "0000011110111100";
		rom(192) <= "0000011101011100";
		rom(193) <= "0000011100011100";
		rom(194) <= "0000011011011100";
		rom(195) <= "0000011010011100";
		rom(196) <= "0000011001011100";
		rom(197) <= "0000011000011100";
		rom(198) <= "0000010111011100";
		rom(199) <= "0000010110011100";
		rom(200) <= "0000010101011100";
		rom(201) <= "0000010100011100";
		rom(202) <= "0000010011011100";
		rom(203) <= "0000010010011100";
		rom(204) <= "0000010001011100";
		rom(205) <= "0000010000011100";
		rom(206) <= "0000001111011100";
		rom(207) <= "0000001110011100";
		rom(208) <= "0000001101101100";
		rom(209) <= "0000001101001100";
		rom(210) <= "0000001100101100";
		rom(211) <= "0000001100001100";
		rom(212) <= "0000001011101100";
		rom(213) <= "0000001011001100";
		rom(214) <= "0000001010101100";
		rom(215) <= "0000001010001100";
		rom(216) <= "0000001001101100";
		rom(217) <= "0000001001001100";
		rom(218) <= "0000001000101100";
		rom(219) <= "0000001000001100";
		rom(220) <= "0000000111101100";
		rom(221) <= "0000000111001100";
		rom(222) <= "0000000110101100";
		rom(223) <= "0000000110001100";
		rom(224) <= "0000000101110100";
		rom(225) <= "0000000101100100";
		rom(226) <= "0000000101010100";
		rom(227) <= "0000000101000100";
		rom(228) <= "0000000100110100";
		rom(229) <= "0000000100100100";
		rom(230) <= "0000000100010100";
		rom(231) <= "0000000100000100";
		rom(232) <= "0000000011110100";
		rom(233) <= "0000000011100100";
		rom(234) <= "0000000011010100";
		rom(235) <= "0000000011000100";
		rom(236) <= "0000000010110100";
		rom(237) <= "0000000010100100";
		rom(238) <= "0000000010010100";
		rom(239) <= "0000000010000100";
		rom(240) <= "0000000001111000";
		rom(241) <= "0000000001110000";
		rom(242) <= "0000000001101000";
		rom(243) <= "0000000001100000";
		rom(244) <= "0000000001011000";
		rom(245) <= "0000000001010000";
		rom(246) <= "0000000001001000";
		rom(247) <= "0000000001000000";
		rom(248) <= "0000000000111000";
		rom(249) <= "0000000000110000";
		rom(250) <= "0000000000101000";
		rom(251) <= "0000000000100000";
		rom(252) <= "0000000000011000";
		rom(253) <= "0000000000010000";
		rom(254) <= "0000000000001000";
		rom(255) <= "0000000000000000";

	end generate;


end RTL;



----------------------------------------------------------------------
--   (C)2005,2006 Copyright J-7SYSTEM Works.  All rights Reserved.  --
----------------------------------------------------------------------
